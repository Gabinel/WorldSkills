��   K�A��*SYST�EM*��V9.3�044 1/9�/2020 A� 	  ����CELL_GRP�_T   � �$'FRAME� $MOU�NT_LOCCC�F_METHOD�  $CPY�_SRC_IDX�_PLATFRM�_OFSCtDI�M_ $BASE{ FSETC���AUX_ORDER   ��XYZ_MAP ��� �LE�NGTH�TTC?H_GP_M~ a �AUTORAIL�_���$$CL�ASS  �S����D��DVERSION�  0��/IRTUAL�-9LOOR qG��DD<x$?������k, � 1 <DwX�< y�����C������	/�� Z�Zm//�/_/�/8�/�/$ �/�/|	?';�$MNU>YA\"�  <� ?/o?'_?�?�?�?�? �?�?�?OOOQO7O IOkO�OO�O�O�O�O�_�O�O_M_�;5N_UM  ��	���92TOOLC?G\ 
Y?-/�_C2  7_�_	o1_o?o%o7o Yo�omo�o�o�o�o�o �o�o;!CqW y������Z�Vy
�Vy