��   �;�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_CPC�_T 4 $�COMMENT �$ENAB�LE  $M�ODJGRP_N�UMKL\  $UFRM\~] _VTX M ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�? �ELAY_T�IMJSPEED�_CTRLKOV�R_LIM? p JD� L��0�UTOO(i��O��&}S. � 8J\TC�u
!����\� �jY0  � ��CHG_SIZ��$AP!�E.�DIS�]$!B�C_+{#s%O#J�
p 	]$Jd#� �&s"��"{#�)�$�'�_S}EEXPAN#�N�iGSTAT�/ DFP_�BASE 5$0K$4!� .6K_V7>H73)&J- � }�\7AXS\UP�CLW�7���
6Jr �< w?�?��?��?�?�// ���&ELEM>/ T �&B�.2NO�G]@%CNH�A�DF#� $DA�TA)
6e0 � PJ�@ 2� 
&P5 ɘ� 1U*n   _VSiSZbRj0jR)(�VyT(�R%S{T_ROBOT�X�S�ARo�U�V$CU�R_��RjSET�U4"	 �bAIS�P_MGN�INP_ASSe#�P B!� `CiH�77`e��.fXc1�CONF�IG_CHK`E_�PO* }dSHRS�T�gM^#/eOTH�ERRBT�j_G]�R�dTv �ku�c
6T1r
0R HLH8�d� 0  lt<N<e'AVRFYhH^tD�5�1� ��W��_A$Rd�TPH/ (G%Q��Q�Q3wBOX/ 8�@F!�F!��G �r{�s"uUI}Ri@  ,��F�pER%@2 {$�p L��_SF��eUIZ}N/ 0 IbF(@�p��Z_�0 _�0wu0  �@�Q7yv	
��~ ��$$CL`  �������Q���Q��VERSI�ON�� � 0��IRT�UAL���' 2� �Q  Q�p���&@>�
m��P�������(������Ғd��Cz  0����A� ��l���������Ɵۯ ���� �2�D�F�h� }�����ԯſ����� 
��.�@�R�d�fϋ� ������п���ώ�� *�<�N�	�rχߖϨ� b��Ͼ�����&�8� ^�\�n߃��߶��� ������"�4�F�X� m�|���������� ���0�B�h�Vx� ����������� ,>Pbw�� �����//( :L�`/��/�� ��/�??$/6/H/ Z/l/�?�/�?�/�/�? �/�?O#O2?D?V?h? jO�?�O�?�?�?�O�O __.O@OROdOvO�O �_�_�O�O�_�O	oo �_<_N_`_r_-o�_�o �_�_�o�_�o)8o Jo\o�o�o�o�2�o �o��o�%�4FX j|��������� ���!�3�B�T�f��� z�������ҏ���� �/�>�P�b�t����� ����Ο������+� =�L�^�p�������� ʯܯ���'�9�H� Z�l�~����ϴ���ؿ ����#�5�G�V�h� zόώ߰�������� ���1�C�R�d�v߈� �߬߮�������	�� -�?���`�r���Q� ����������; M\�n���������� V����"7IX j|������ ��/E/W/fx ���/��/��/ ?,/A?S?b/t/�/�/ �/�?�/�?�/?O(? =OOOaOp?�?�?:O�O �?�O�? OO'_6OK_ ]_lO~O�O�O�O�_�O �_�O_#o2_GoYoko z_�_�_�_�o�_�o�_ 
o@o1 Ugvo�o �o�o�o�o�� -�<Q�c����� �u�����Ώ8� *�_�q�������ʏȏ�ڋ�$DCSS_CSC 2����Q � P����:�܉d 
�k�.���R���v�ׯ ����Я1���U�� y�<���`���ӿ���� ���޿?��c�u�8� ��\Ͻπ��Ϥ���� ��;���_�"߃�Fߧ� j߷��ߠ����%��� I��m�0���f����������GRP ;2�� ����	ҟS�>�w�b����� ����������= (aL�p��� ��� K6 oZ�~���� ��/5/ /Y/D/}/ h/�/�/�/�/�/�/? �/
?C?.?g?R?�?�? �?z?�?�?�?�?O-O OQO<OuO�O�OdO�O �O�O�O_�O_;_&_ __q_�_N_�_�_�_�_��_�_�_%ooIo��_�GSTAT 2���%��< ��2�R�4���!?�  �a5�����fRߵ���ɘa��Q%�� D4��C���U��8`<�e�q��?x�Y����ƫ�����b�`>�`4��Z����C�8�����e>Gҿ��}?IDT>�=��C�!��3��iBPU���V��C��� y��C.>ّ�2?f:F�x��X�`��=��>�Y>��_��>����A������D"�k y���Q����]��IJ5>Y?�dtϿfRǵa�lV>�}�`�D�bVxz�}��L�q?�p5�()�p�5A�{뿙`4�Q&� �o�o�o y��<�N��� 0�z���f���Љ�i �-i��+k y �.�� &�H�v�\�~������� �ȟڟ��*���Z�l� ��x���|���د��� .��B��J�0�B�d� ��x���ȿ������� ���F�H��Ϻ�t�����Ϫ�����͵����?�6<��R����t��j���P4�����5@�K��C�"D)����m<rE�?����b���1�~ɯ�qмm��a@���C���m��Mq�YR?���� gʿ�ٿYe������ó`�C�� y��Q�>��� ?r��;�q�<rDN�����eњ��r�p������Ǹ����Cw�ް�ڌ�-��}���:�e�� ��p��pK&����@�MCĿڑDB�� y<�p]�?�)<��MJ���<pK�9��/5��}�I�0�O�F�(�:� L����������� ��� �V�h��Pϒ�dϪ� ����������F ,^|bt��j� �8��<N(r �z������� ��,//4/b/H/Z/ |/�/�/�/�/�/�"? T?X?j?D?�?�?z? ���P�b�t߆ߘߪ� ����������(�:� L�^�p��O�?�?�?�? t_�_|?�_�_�_�_�_ o��/.o ?FodoJo \o~o�o�o�o�o�o�o �o2`?�� �_����� �o dJ�xB�d���x��� ȏ��Џ������F� ,�N�|�b�(������ �����*�<��4_F_ �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O _~�`�r�����"� �.�X�2�DώϠ�:� ���Ϝ��� ������ H�.�P�~�dߖߴߚ� �����ߢ�,�>�p�*� t��`���� ��� ��� �.��6�d�J� l��������������� ����Z��F�� |���п⿈��� ����Я�����*� <�N�`�r�������/ � ��/�/��/ �/�/�/*?<?��$f? 8~?�?�?�?�?�?�? �?O O2OPO6OHOjO �O>�O�O?�O_"_ �OF_X_N?�O�_�Oz_ �_�_�_�_ o�_o6o o.oPo~odo�o�o�o `_�o(_�o,>b tNl/~/$6HZ l~������ �/ /2/D/���� �VH�Z�Pf���j� |�Ɵ؟r_�o��o� 8��0�R���f����� ��ί�ү��4��o d�v���b�������� ���8��L��8�f� L�nϜςϤ��ϸ��� ��� �"�P�6����� Ŀ~����ߴ������ �������� ,�>�P�b�t������� ��Ώ��R�4�F�X��� ������,b t�\ߞp߶�� ��$R8j �n���v� // D�H/Z/4/~/�/� ��/��/�/?�/
? 8??@?n?T?f?�?�? �?�?�?�?�/.O`/O dOvOPO�O�O�O���� \�n��������� �����"�4�F�X�j� |��_�O�O�O�O�o�o �O�o�o�o�o�o�/ �?:ORpVh� ������$�
� �>�l�O�����o�� ���Џ�,�"p�V� ��N�p�������ԟ�� ܟ
���$�R�8�Z� ��n�4�ʯ���� ����6�H�V��$DC�SS_JPC 2�@�Q �( DMP���� ����P��ۿ����� ���Y�(�g�Lϡ� p��ϔ��ϸ����1�  ��g�6�H�Z߯�~� �ߢ��������?��  �u�D�V�h����� �����)���M��.� p���d�v��������� ��7[*N �r�����! �/i8�\� ������//� /"/w/F/�/j/�/�/ �/�/?�/�/=??? 0?�?T?�?x?�?�?�? �?O�?�?8O]O,O>O �ObOtO�O�O�O�O�O #_�OG__k_:_L_�_ p_�_�_�_�_�_��h�Sq�u�L�_Uooyo��dDo�oho�o�o �o�o�o1�oU y@Rd���� ���?��c�*��� N���r�����󏺏̏ ޏ��M��q�8���\� ����ݟ���ȟ%�� ���Y��F���j�ǯ ��믲��֯3���W� �e�B���f�x����� ������A��e�,� ��Pϭ�t��ϘϪϼ� �+���O��s�:ߗ� ^߻߂��ߦ����� ��K��$�6�H��l� ���������5��� Y� �}�D�V�h����� ��������C
g .�R�v��� ����Qu< �`����/��&dMODEL 2�3kx��
� <�c (  �z(�/g/y/ �/�/�/�/�/�/�/D? ?-?z?Q?c?u?�?�? �?�?�?�?.OOO)O ;OMO_O�_�OY/�O�O _�O�O<__%_7_�_ [_m_�_�_�_�_�_�_ �_8oo!onoEoWo�o {o�o�o�o�o�o�O�O �O�o|�oew� �����0��� +�=�O�a�������� ��͏ߏ���b�9� K���3Es����m� ۟����#�p�G�Y� ��}�������ůׯ$� ���Z�1�C�U�g�y� ��ؿ����ϩ���� ��h��Q�cϰχϙ� �Ͻ��������d� ;�Mߚ�q߃��ߧ߹� ������N�%�7�� �1�C�q��Y����� &����\�3�E�W�i� {������������� /A�ew� ��������� �=O�s��� ����/P/'/9/ �/]/o/�/�/�/�/? �/�/:??#?5?�? /]?o?�?�?�?O�? �?HOO1OCO�OgOyO �O�O�O�O�O�O�OD_ _-_z_Q_c_�_�_�_ �_�?
o�?�_�_Ro)o ;o�o_oqo�o�o�o�o �o�o<%7I [m������ ���!��_��oI� [�ȏ������Տ��� ��/�|�S�e����� ������џ�0��� f�=�O�a�s�����m� ������ѯ>��'�t� K�]�o��������ɿ ۿ(����#�p�G�Y� ��}Ϗ��ϳ�����$� �������5�Gߴ� /ߝ߯�������2�	� �h�?�Q�c�u��� ����������)� ;�M���q�����k�}� ����*��%7I [������ ��\3E�i {����/�� F/����!/3/�//�/ �/�/�/�/?�/?T? +?=?O?�?s?�?�?�? �?O�?�?OPO'O9O �O]OoO�OW/i/{/�O �O�O�O_^_5_G_�_ k_}_�_�_�_�_o�_ �_Hoo1oCoUogoyo �o�o�o�o�o�o�o�O V�O1u�� ��
�����)� ;���_�q��������� ˏݏ�<��%�r�I��[�m����$DCS�S_PSTAT ����ӑ�Q    ��� � (��+��O���t� r�Ԑ�������������ӕ௎�կ��ĔSETUP �	әBȖ��� ��8�R�ͬs�b����������T1SC 2i
+�����Cz�������صCP R-�D�DLj� |�>�ϲ��ϓ����� ���0�B�T�#�xߊ� Yߛ����ߡ����� ��>�P�b�1���� y��������(��� L�^�p�?��������� ��������$6Z l~��Vϫ�D� ��);Mq ��d����/ /�7/I/[/*//�/ �/r/�/�/�/�/?!? �/?W?i?8?�?�?�? �?�?�?�?�?O/OAO OeOwOFO�O�O�O� �O�O_�O+_=_O__ s_�_�_f_�_�_�_�_ oo�_9oKo]o,o�o �o�oto�o�o�o�o #�oGYk:�� �������1�  ��g�y�H������� �����	��O-�?�Q� ؏u�����h���ϟ�� ����;�M�_�.� ������v�˯ݯ���� �%���I�[�m�<��� ������ٿ���̿!� 3��W�i�{�Jϟϱ� �ϒ��������/�A� S�"�w߉��j߿��� ��������=�O�a� 0����x������ ��'���K�]�o�>� ���������������� #5Yk}L� ������1 Cgy�Z߯� �Z�	//�?/Q/ c/2/�/�/h/z/�/�/ �/??)?�/M?_?q? @?�?�?�?�?�?�?�? O%O7OO[OmOONO �O�O�O�O�O�O�O�O 3_E__i_{_�_\_�_ �_�_��_oo�_Ao Soeo4o�o�ojo�o�o �o�o+�oOa sB��x��� ��'�9��]�o��� P�����ɏ�����Ώ #�5�G��k�}���^� ��şן�������_ C�U�ܟ6�����l��� ӯ寴�	��-���Q� c�u�D�����z�Ͽ� �¿�)�;�
�_�q� ��RϧϹψϚ���� ��%�7�I��m�ߑ� `ߵ����ߨ�������3�E�W�&��$DC�SS_TCPMA�P  ������Q @� .�.�.�T.���.�.�.�U.�	.�
.�.�U.�.�.�/�W  .�.�.�U.�.�.�.�.�.�.�.��.�.�.�.� �.�!.�".�#.�$�.�%.�&.�'.�(�.�).�*.�+.�,�.�-.�..�/.�0�.�1.�2.�3.�4�.�5.�6.�7.�8�.�9.�:.�;.�<�.�=.�>.�?.�@�u�UIRO 2.��������� ������,>P bt�������-���-��Q cu������ �//)/;/M/_/q/ �/�/2�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O�/ 3O�/WOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_&O�_q�UIZN 2��	 ����� oo $o*��_Rodovo9o�o �o�o�o�o�o�o* <Nr��Y� �����&�8�� \�n�=�������ȏ�� ����ߏ4�F�X�� |�����o�ğ֟蟫� ��0���T�f�x�;� M������������_~x�UFRM R�����81�^�p� /����ʿܿ�� � ��6�H�#�l�~�Y� �ϴϏ��������� � 2�I�V�h�ߌߞ�y� ���߯���
���.�@� �d�v�Q����� �������*�A�N�`� �����q��������� ��8J%n� [������ "9�FX�|�i �����/�0/ B//f/x/S/�/�/�/ �/�/�/??1(?P? b?=?�?�?s?�?�?�? �?O�?(O:OO^OpO KO�O�O�O�O�O�O _ _)?;?H_Z_�O~_�_ k_�_�_�_�_�_�_ o 2ooVohoCo�o�oyo �o�o�o�o
3_@ R�ov�c��� ����*��;�`� r�M�������̏ޏ�� ��+8�J��n��� [�������ǟ���ٟ "�4��X�j�E����� {�į֯������