��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ��!PCOUPLE�,   $�!P=PV1CES0�!H�1�!"PR0�2	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U}4 Q �ARG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W�1�W 6P!SBN�_CF�!�0�$!J� ; 
2�1_�CMNT�$F�LAGS]�CH�E"$Nb_OP�T�2k�(CEL�LSETUP 7 `�0HO�0 �PRZ1%{cMAC{RO�bREPR�hD0D+t@��b{�e[HM MN�B
1^ UTOB U��0 9DoEVIC4STI�0��� P@13��`B�Qdf"VAL�#IS�P_UNI�#p_�DOv7IyFR_F�@K%D13�;A�c�C_WA?t�a�z�OFF_@N�DEL�xLF0q�A�q�r?q�p�C?�`�A�E�C#�s�A�TB�t�D�MO<� �sE � [�M�s��2�REV��BILF��XI�� %�R  �� OD}`j��$NO`M�!b�x�/�"u�� ��������@Dd� p E RD_�Eb��$FSS�B�&W`KBD_S�E2uAG� G�2B "_��B�� V�tp:5`ׁQC  ��a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR�� BIGALLOW� (KD2�2�@VAR5�d!�A�B �BL[@S �C ,KJqM�H`S�p�Z@M_O]z��w�CFd X�0�GR@��M�N�FLI���;@UI�RE�84�"� SW�IT=$/0_No`S��"CFd0M�{ �#PEED��@!�%`���p3`J3t	V�&$E�..p`|L��ELBOF�  �m��m�p/0��C	P�� F�B����1x��r@1J1E_y_T>!Բ�`��gt���G� �0WARNMxp�d�%`�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�M�� R�r$OR�I�.&ӧRT�S�Fg CHGV0I��p�T��PA�I�{�T�!��� � �#@a����HDR�B��2�BJP; �C��3�4�U5�6�7�8��9�4��x@�2 ]@� TRQ��$%fh��ր����_U����B�COc <� ����Ȩ3�2�ЯLLECM�-�MULTIV4�"$��A|
2q�CHILD>��
1D��z@T_1b � 4� STY 2�b4�=@�)24�p���?�� |9$��T�A�I`�E���eTO���E��EXT���ᗑ�B��2G2�0>��@���1b.'��B ��A�K�  �"K�/% �a��R���?sA�>�O�A!M��;A�֗�M�� 	�  =�I�" L�0[�� R�z�pA��$JOBB�x�����TRIGI�# dӀ����R��-'r��A�ҧ��_M���b$ tӀFL�6�BNG�A��TBA� ϑ�!��
/1�@À�0���R0�P/pX ����%�|���Bq@W�
2JW�_)RH�CZJZ�_*zJ?�D/5C�	͠ӧ��@���Rd&�������ȯ�qG|Өg@NHANC��$LG/��a2qӐ� ـ��A�p� ���a�R��>$x��?#D�B�?#RA�c?#A�Zt@�(.�����`F3CT����_F࠳`&�SM��!I�+lA �%` �` ���$/��/����[�a��M`�0\��`��أHK��CAEs@͐�!�"W���N� SbXYZWȝ`�"����6	��j�I��'  E. II��2�(p�STD_C�t�1Q]��USTڒU�)#�0U[�%?I-O1��� _Up�q��* \��=�#AO�Rzs8Bp;�]��`O,6  RSY�G�0�q ^EUp��H`G�� ��?��@PXWORK��+@�$SKPa_�p��A�TR�p , �=�`����Z m�OD3��a �_C"�;b�C� �GPAL:c�a�tőS�D�W�3Bb����P���P� @�!�-�B APR��

�qDJa3��. /��u�������LuY/$�_����0�_��/�PC�1�_����~�EG�]� �2�_���AF�.��R3�H $C��7.$L8c/$uSނ�z IkINE�WA_D1%�ROyp��ŀ����q�c7 t@�fP�A���RETUR�N�b�MMR"U���I�CRg`EWM�@�SIGNZ�A� ���e� 0{$P'�1$P� &m�2p�p'tm�+pD�@ �'�bdNa|)r�GO_AW ���@ؑB1TPCYSd�(�CYI�4��B�`1w�qu��t2�z2�vN�}��E}s�DEVIs` 5� P $��RB���I�wPk��IG_BY���"�T7Q��tHNDG�Q6� H4��1�w��$DSBLC��o��v�g@��j}sL��70O�f@]���FB���FEra8�ׂ�t}s��
�8> i�T1?���MCS���fD �ւ
[2H� W��EE����%F���I�q����9� T�p��x�NK_QN:�����U��L�wKHA�vZ' ~�2�p���v�q7: �='MDLn���9�ጂ ٱh����!e����J��~�+����,�N�D����3��ՒG��AqSLAd�7;;  ��INP��"�`����}q_ �4<�0�6`C� NU��+  D�LקRR��SSH!�7=M��q���ܢӢ����sP���>P +$ٰ�٢��^��X^�Y�FI B\�@�Ă��'A	'AWl�N��NTV��]�V~�.X�SKI�#T����a�ۺ�T1J�3:3_�P�SAFN����_SV�EXCL�U��N@�DV@L���@�Y����S�HI�_V
0\2PPLYPRo�HIM�T�n��_MLX��pVR�FY_�Cl�M��I3OC�UC_� �d���O�q�LS�0�M2FT4Q������@P�E$�t��A��CNFK66եu�8�pm�4ACHD�o�ؕ����AFC CPDlV�TQ����_��g ?`�@TA�@��0L@ �Q��N���]� @����T��T! S����te@{R�A DO�� w23���!n��	_1�#�H!� b�� �΀K��B�2��MA�RGI�$����A���{s_SGNE�C;
$�`�a^aR0 ��3��@ B��B��ANNUN�P?����uCN@�`%0��`��� ���BEFc@]I�RD @Q�F���4OT�`�sFTӠHR,Q��CQ0�M��N�I|RE�����A�W���DAY=CLOCAD�t;T|�<S5CQ�j�EFF_AX�I��F`1QO3O���S�@_RTRQ�E�G����0RQ
�2Evp ��ꐁF�0f�R0 �t��AMP�E<� H 0�`œ^��`Ds�DU�`��v�BCAr� I?��`N ErIDLE_PWRI\V!n0�V�wV_[ ꐅ ��DIAG�5J�o 1$V�`SE�3TQl�e��P�l�^E_��Y�VE6� �0SWH�q (� �b�Gn�3OHxPPHZ�IRAl�B�@�[� �a�b�1�w3�O  � ��v��I�0 ��pRQDW�MS-�%AX{6Y�LIFE�@�&�MQy�NH!Q%��F#�C����CB0�mpNr$�Y @�aFLAl�f��OV0]&HE��>l�SUPPO�@L1�y��@_�$��!_�X83�$gq�'Z�*W��*B1�'T�#`�k2XYZáY�Y2D8CY`T@�`N����f� �C�I2��� C�TA�K `�pCACH�ӫ�3�����I��bNӰUFFI� \��@��;T��r<S6CQ�MSW�5�L 8	�KEYI7MAG�cTMLa���*Ax�&E���B;�OC�VIER-aM ���BGL����y�?��I�"`�П4N�6:�ST�!�BP��D,P�D��D��@EMAI䐔a����s�/FAUL|RObB�c��� spUʰ�`��T�'`E�P< $dS�S[ � ITw��BUF�7y��7�tN�[�LSUB1T�C�x�o�R�tRSAV |U>R'c2�\�WT����P�T�*`Sn�_01PbU���YOT�bK�
�P��M��d���W#AX��2��X1P�ְS_GH#
��YN�_���Q <Q�D���0���M�*� T�F�`|�\�{DI��EDT_P$ɰ:�R��b�GRQM�&��Jq�a�1׀��F�s� S (�SVqpB��4�_���a~��T� �@����B�SC_R]1IAK>B'r��$t��R"A8#u�H�aDSP:FrP�lyIM|Sas�qz��a� U>w� <1%sM�@IP��s��0�`tTHb0ЃTr��T�`asHS�cCsBSCʴq0� V�����S�_D��CONVE�G���b0^v1P	FHy�dCs�`&a?A�SC���sMER|g��aFBCMPg�v�`ET[� UB�FU� DU%P�D�:12�CDWy�p�PD�CpR��6�:�V� ��� ���P���C"�����w�����|`��WH *�LƠ�Cc�W����Y� 賂��р�q�|�P��A��7}�8}��9}�H ���1��1���1��1��1ʚ1�ך1�1�2��2T����2��2��2��U2ʚ2ך2�2�3��3��3����3���3��3ʚ3ך3��3�4�����O�EXT[�X[b �H``t&``z�k`˷$���0FDR�YTPV��RK"	�\�K"REM*F��N]"OVM:s/�A8�oTROV8�DT�P6X�MXg�IN8ɉ �W��INDv�H2
�ȕ`K ^`G1a�a�Ȉ@Q%7Da�RI�V��u"]"GEAR�:qIO.K(�H4N �`���,(�F@� I3Z_MCM<0K!��r� UT���Z ,��TQ? b�y@\t�G?t�E  |�PA>Q����[p�5Pa� RI�E@�>SETUP2_ g\ �@=STD	p<TT�������Ֆ1�>RBACUb] T(��>R�d)�j%C�E��0��IFI��0���i�{�4�PTT�AF�LUI�D^ �� gHPUR�gQ�"@�r�a�4P+ I�u$��Sd�?x���J�`CO�P�SVR�T��N�x$SHO8* ��CASS��Q8w%�pٴBG_%��3����F�ORC�B��o�DAkTA��_�BFU_�	1�bb�2�a�an�b0���` |��NAVN	`������$��S�Bu#$VIS�I���2SC	dSE������V��O��$&�BK�� ���$PO��I���FMR2��a ��	��` #��&�8�O� �(�_����+IT_^�ۄ)M������DGCLF�DG�DY�LD����5�Y&��Q$��M됇Cb�N@{	 T�F9S�P�Dc P��W|�cK $EX_W�nW1%`]��"X3��5��G+�d� ���SWeUO>�DEBUG���-�GR��;@U�B�KU��O1R� _ PO_ )���t��M��LOOc>!SM� E�R�����u _E e �>@��0TERM�`%fi%M_M�O�RI�ae gi%��S#M_�`>Re hi%X��V�(ii%����UP\Bj� -����e��w#� f���G�*ELTOr�A�bF�FIG�2��a_���Ў$�$g$wUFR�b$�01R0օ� OT_7F��TA�p q3NST��`PAT�q�0�2P'THJ�ԀE�@�c3ART�P'58�Q�B�aREL�:�aSHFT�r�a�1�8E_��R��у�& � 	$�'@i�
����sN@bSHI�0�Uy�~��$PAYLO�p �Oaq�����1����pERV��XA��H ��m7�`�2%�P�E3��P�RC���ASY1M�a��aWJ07�����E�ӷ1�I��ׁU�T�`Oa�5�F�5P��su@J�7FOR�`MF 
�O!k]���5&�0L0��`HOL ;l �s2T����OC1!E�$OP��qn���#$�����$��P�R^��aOU��3e��R�5e�X�1 ��e$PWR��IMe�BR_�S�4�� �3�aUD��k�Q�d]m��$H�e!�`�ADDR˶HR!GP�2�a�a�a��R��.[�n H��S����%��e3��e���e��S�E��z�HS�MNu�o���P��q��0OL�s߰`xڵ�I ACRO��<&1��ND_C�s�x�AfdK�ROUP�B�R_�В� �Q1|� =�s���y%��y-��x@���y���y>�=A��<Ҁ�AVED�w-���u�P(qp $_��P_D�� ��'r�PRM_�� �HTTP_��H[�q (ÀOB�J��b �$˶L�E~3�\�r � Q���ྰ_��TE#�ԂS�PIC��KRL~PiHITCOU�!��L���PԂ���0���PR��PSSB�{��JQUERY_F�LAvs�@_WEBwSOC���HW��#1��s�`<PIN'CPU(���O��� g�����d��t��O��C�IOLN�t� 8��R��$�SL!$INP7UT_U!$`���P M֐SL.���u���2�.���C��B��IOa�F�_AS=v�$!L+ਇ+�A��bb�41�����Z@HY�ʷ�����!e�UOP:w `v�ϡ˶�� ��������"`PIC`����� �	�sQIP�_ME��v�x X�v�IP�`(�R�_N�p�d���Rʳp�ױQrSP �z�C��BG(�OG���M��Av�y l�@CTiApB��AL TI�`3UfP_ ۵�0PSڶBU_ ID� 
�L �� `šQ����0�z)����ϴ�N�N�_ O��IRCA�_CNf� { ��Ɖ-�CYpEA��������IC����tpR�=QDAYy_
��NTVA������!��5����SCAj@��CL�
����
���v�|5�VĬ2,b�l�N_�PCV�n�
���w�})�T��S�р���
��e���T� ?2| �� ��v�~��֣�ذLA�B1��_ ��UNIrX��ӑ ITY����e�!IR� ��<�)���R_URLn���$A;qEN ����s`vsTeqT_�U���J��X�M�$���E�ᒐR�祪�� A�,���J�H���FLy��= 
|���
�UJR|U� ���F�6G���K7��D>�$J7,�s��J8*�7���$3�E�7��&�8\�)�oAPHIQ4�zy�DkJ7J8Rޒ�L_KE'� o �K͐LMX�� � <U�XR�i�����WATCH�_VAZqu@AំF'IEL`��cyԐ��&:� � u1VbwPFCTX�j���LGE��� �!��LG_SIZ�΄�[8Zm�ZFDeIYp1!gX b ZW �S`�8� m��� �b ��A�:0_i0_CMc3#�*'FQ1KW rd(V(Bb�po pm�p� |I�o�1 pb pW RyS��0  (r SLN�R�۠�DE6E3����c��i���PL#�DAU"%EAq�͐�T8"�. GH�R�!y�BO�O�a�� C��F�ITV�l$A0��sRE���(SCRX�����D&�ǒ�qMARGI�Sp�,�����T�"�y�S��x�Wp�$y�$��JGM7�MNCHt�y�FNĤ�6K@7r�>9UF�L87@L8FWDL8H]L�9STPL:VL8�"�L8s L8RS�9HOPh;��C9D�3R��}P�'IUh�`4�'��5$ ��S2G09�pPOWG�:�%�3,64��vN9EX��TUI>5I� �ӌ�����C3�C<0'�,�o:��&��@�!NaqvcANAy��Q�AI]�gt7���DCS���cRS�c*RROXXOdWS�ÂRroXS{X�(IGNp �
Ђ=10 ��[TDEmV�7LL��
Z!�*�C �	 8�Tr�$f/蛒��m��3A�a�	 W�萦�ZOqs�S1Je2Je3Ja���ASPC G� �ƋG`-T� �%��Q�T�r@�&E�V�fST�R9 YBr~�a �$E�fC�k�g��f	v(e� B� L����� �� u�xs뀔�g�q�jt����"�#_ � �[��w�#Ӡ �s �{MC�� ����CLDP᠜�TR�QLI ���y�tFAL���rQ��s5�D���w~�LD�u�t�uO�RG���1�RESERV��M���M��Œ�s��� �� 	�u�5�t�uSVH��p��	1�����RCLMC��M�_��ωА����MDBG�h�I����$DE?BUGMAS�������U�$T8P��E�F�d�C�MFR�QҤ� � ~K	HRS_RU��bq��A��$EFR3EQ6u!$0YOVER�k��f��PU1EFI�!%Gq�� �aMY�z�ǐ \����E�$9U�`��?��
�SPSI`��	��CA ���ʲ�σUY�%��?( 	�MIS�C�� d��aR5Q��	��TB� �c ���A��AX����𑧪�EXCESHg�W!d�M�H�9�au����Qd�SC�`� � H�х�_�����������נK�E��+�� &�B_^, FLICBtB� �QUIRE CMO�t�O������MuLdpMD� �p�{!��5b���n�M#ND!��I�����L �D;
$INAsUT�!
$RSM�ȧPN�b�C�j`��PSTLH� �4U�LOC�fRI�"��eEX��ANG�.R.�~p� A]��bq��� ���MF0 ����icr�@mu����$�SUPiu�qFX��IGG! � ���cs��#cs
F ct��ޒ�b5��`E��`�T�5�tC��g�TI���C`r�� M����� t��MD���) ��XP��ԁ��H��.���DIAa��Ӻ�W��!��0af���D@#)�a�O�㥀��� �CUp V	���.����O�!_��ᜃ �{`�c����	�� |�P|��0� ���P{�KEB��e-�$B��o�=pND2xւ����2_TXlt�XTRAXS����&��LO: ����&}�M���C�.��&�`�RR2h���� -�!A�� d$CALI����GFQj�2F`RI�Nbn�<$Rx�S�W0ۄ���ABC��D_J��{�T���_J3��
��1S�P, �T�P����3P��H�9pT�#J�h3n���O�QIM�M�CSKP�zb7$?SbJ+�M�Qb�py����_AZ���/�EL�Q.ցO�CMP��N�� R1TE�� �1�0 �F��1��@ Z�SMG�0����JGΊpSCLʠ��SPH_�PM��f��T�=u�RTER��n�IPk�_EP�q�`aA� �cM��DI��Q23UdDF � ���LW�VE�L�qINxr�@�_�BLXP.��Y/�J`��'$X IN���]�C�9%�"T�7":6p_T� �F%a"���^$��k)�j`�DHʠ��\�9`�$Vw��_�A$�=����&A$���נR6�]�H �$BEL� m���_ACCE� x	8�0IRC_��q�@�NT��c�$PSʠ�rL� ��M4�s9 .7��GP/6 ��9�7$3�73S2T�͡_Ga�"�0�1��8�n1_MG}�DD�1���FW�p��3�5�$32�8DEKPP�ABN[7ROgEE�2KaBO�p�Ka���1�$USE�_v�SP��CTR�TY4@� �� <qYNg�A�@�FR �ѢA!M:�N�=R�0O�v1�DINC(��B�4p���GY��ENC��L��.�K12��H0I�N�bIS28U��ON�T�%NT23_���fSLO���|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1���M�PERCH  �S��� �W���Sl� �R��l����E�0�0PAS2EeL�DP7��ONUЉZ�f�VTRK�RqAY"�?c� �aS2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gB�T�DUX �2S_BCKLSH_CS2 Fu:��V���C-�esR�oz�A�CLALM�JT@��`� �uCHK�e ����GLRTY@pн�8T��5���_��N�T_UM3��vC3�p�1Z���LMT���_LG��%���0�E *�K�=�)�@5F�@8 09�Nb��)hPC�Q)h�HТ��5�uCMC����0�7CN_��N����;SF�!iV �B��.W���S2/�Ĉ7CAT�~SH�Å� �4 V�q/q/V�T1���0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e�0�R� @B�_Wu�d��!a��#`��#`�I*h�Iv�I�#F��S��:��I�0VC00��֢1ܮ�0��JRKܬ!��<�KDBXMt�<�M��_DL�!_bGRV�g�`��#`��#A�H_p%�?��0��COS��� ��LN#���ߥŴ � ��=������꼰�b<�Z���VA�MYǱ�:ȧ��᯻[�THE{T0�UNK23�#؅��#ȰCB��CB�#Cz�AS�ѯ�0���#����SB�#��N��GTSkZAC�������&���$DU�phg6�j��E��%Q%a_��x�NE
hs1K�t�� y�A}Ŧկ׍������LPH����^U��S ߥ����������!�(�(Ʀ�V��V�غ ���V��V��V
�V��V&�V4�VB�H���������d�����H�
�H�H&�H4�H*B�O��O��Os���UO��O��O
�O�UO&�O4�O(�F����	���SPBALANCE_J��6LE��H_}�S�P>!۶^�^��PFULCb�q����K*1�UTOy_�p�uT1T2�	
22N�q2VP�M@�a� i�Z23	qTu`�O� 1Q�INSE9G2�QREV�P�GQDIF�ep)1�lU�"1�SPOBK�qj�w2,�VP�qI�?LCHWAR4B�B�AB��u$ME�CH��J��A��vAX�aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ֯@�C1_ɒT �� x $W�EIGH�@�`$ȹ�\#��I�A�PIF�vA�0LAG�B��S��B:�BBIL�%O1D�`�Ps"ST0s"P:�pt �� N�C!
L �P 
P2�Aɑ�  2��Tx&DEKBU�#L|0�"5�OMMY9C59N���$4�`$D|1 a�$0ېl� �_ �DO_:0AK!� <_ �&� �q�A���B�"� NJS�8_ԍP�@��"O�p _�� %�T7P�?Q�TL4F0TI�CK�#�T1N0%�3=p�0N�P� u3�PR\p�A��5��5U0_PROMP�CE��? $IR"��Ap�p8BX`wBMAIF�h�A�BQE_� OC�X�a�@RU�COD��#FU�@�&ID_��P�E82B> G_SwUFF�� �#4�AXA�2DO�7/�5� �6GR�#��D C�D��E��E-��D�U4� �_ H_F�I�!9GSORDf�! R 236s��HR�AN0$ZDT�E=!� X5�4 =*WL_NA�1�0|�R�5DEF_I�X �RF�T�5�"�6�$�60�S�5�UFISm�#� m1|��40c�3�T6�"44􁆂�"D� ?r�fd�#D�O@ l2LOCKE���C�?O0G2a�B�@UM�E�R �D�S�D�U�D>b�B�c �E�S�Dd�B�&2v2a �C�ʑ�E�R�E�S�C9wwu�H�0P} d�0�,a��F0W�h�u�c�=!TE�qY4�� �!LOMB_t�r�w0s"VIS��WITYs"AۑO�#A_FRI��~#SI,a�n�R�07���07�3�#s"W�W��Q��%�_���AEAS{#�B��|�x`TWB8�45�55�6|#�ORMULA_I�G�W� h� 
>75COEFF_O�1&)��1���Go�{#S� 52CaA� :?L3�!GRm�� � � $h�`�v2X�0TM�g����e�2�c��3ER�IT�d�T� �  ��LL�Dp`S��_3SVkd��$�v� q�.���� � ���SETU,cMEA�G@�@Πt �!HRL �� � (�   0��l��l��aw��R��0�a�a}d]� d��B��Ay`Gax`賫[Ѐk@RECt[Qq��!SK_A �y�� P_!1_USER����8*���VEL�����-�!��IzPB��MT�1CFG���O  �0]O��NOREJ �0l����[�� 4 pe���"�XYZ<S�B� 3:!��_ERRK!� U ѐ�1�@Ac�Ȱ�!�>�B0BUFINDX���ñMORy�� H_ CUȱ�1���dAyQ?�I>Q�$ +�a�����ñ\�G{�� ?� $SI�h��@2	�VOv�q�- �OBJE| w�ADcJUF2yĈ�AY��4���D��OUKP�����AMR=�T���-���X2DIR�����Xf�1  DY�Nt�0�-�T� ��R���0� ���OPW�OR�� �,>B0SYSBU�����SOPo���z�U�y�XP�`K���PA`�q������OP�@U���}�"1��/IMAG۱_ ��f�"IM.���IN�������RGOVRD"ё�	���P����  �>gplcC��L�`B�Ű?l�PMC_E(�P�1N��Mr�1b212��"�SL| ���� �R OVSuL=S�rDEX\aD`��2�:�_"� ��P#���P������2�C �P>���^#�_ZERl���:���� @��:��MO�@RIy��
[�`g@e���s�Q�PL����  $FR+EEY�EU��Z*��L����T�� �ATUSk�,1C_T�����B�������p�Vc1��P��� !Dc1�к���LQ��`��MQ��ۡL�XE�� x�5IP�W�` ���UP��H`&aPX�;@��43����PGY��g�$SUB���q���JMPWAIT~ ���LOW���1w�� CVF_A�0���R�Z��CC �R�$��28IGNR_{PL��DBTB� P*a�BW@.t��U�0-IG��!@I��TNLN,�R�Bѡb�N!@��PE�ED~ ��HADO!W� ��t���E�������PSPD��� L_ A�нP��Æ	#UNq � �R�P (�LYwPa��~N �PH_PK����b�RETRIE��x���)�PS D@;FI��� ���V ރ$ 2�d�DB�GLV<LOGS�IZz�baKTU����$D��_TXV�EM�Cڡ)�� ��-R�#�r��CHEsCKz��	�PL�J��ϰq)�L��.��NPA�`TJ"��J��*0P����
�AR�"�BC =Sa��qO�@����ATTS� u䡳&� w�^a�3-#cUX^�4�QPL�@�Z�� $d��qSWOITCH�h�W��{AS�����4�LLB��� /$BA�Dvc���BAMi��6I��F(@J5��N�UB6[F>
A_KNOWK3qB"�U��AD+Hc� �D��IPAYLOAq�9p�C_���Gr�*�GZ�CLqAj��P�LCL_6� !�4��BOA?�T7�
VFYCӐ�Jp��D
�I�HRՐ�G�T�B��6�J(�zQ_Jt�A �B�AND�����T�BQP���PL~@AL_ ��0� =�TAe��pC��D:�CE���J3�P�V�� T�PDCK�^�)b��COM�_AgLPH�ScBE<�߁�_�\�X�x\�� � ���OD�_1�J2�DDM�A�R<�h�e�f�cQ�TWIA4�i5�i6��MOM(��c�c�c�c4�cV�B� AD�cv��cv�cPUBP�R �d<u�c<u�bf�2����� L$PI $��pc��G�y��I*�yI�{I�{I�s�`@�A���v��v�J��b��a��HIG �3���0���5 �0�f�?�5N�5�SAMPD Ƣ�0�p���;@�S �� с6���1���� �� �`���`1�K�P��`�d�P�H��IN1� �P��8�T�/��:�z�xQ�z���GAMM&��S��$GET������D^d>�
$N�PIBR��I��$HI��_���1��E=��A�9�*�LW�W�N�9�{�*��Zb���QCdCH�K0�j�ݠnI_ ��M�JļRoh�Q ���sJ�-v��S {�$�X 1�N�}I�RCH_Dx!�$RN���^�L�E��i�p�Zh8�ž�MSWFL/Mn�PSCR�75��� ��3�"Ķ�6��``��ع���4SV���P'������G�RO�g�S_SA�=AH�=ńNO^`C i�_d=��no�O�O �x�ʚ��p�B�u�ȐcDO�A��!�ں �*�t�:�Z1f�;�7�����CFMmu� � �YL�snQ ��� ���"��<s�	�����nQ૰<N3M_Wl�����\p��(�o�MC��P���Q����rhpM.�pr� ��!ȅ�$�WM��ANGL�!�AM�6dK�=d@K�DdK��TT7�Nk@P��3�#�PXC OEc¼QZ��hp	nt� -���OM���� �ϣϵ����`� c�Z0tes^a_�2� |a �J��i���c���cJ���j�����jA� (�z����0�@{��P�1�PMON_�QU�� � 8�60QCOU��Q�THxHO��B H�YS�0ESPBB U�E- 3�f0O�4� � c P�^�RU�N_TO���0O��� P�@���INDE�#_PG�RA���0��2��N�E_NO��ITxf��o INFO���a"������1O�I� (*�SLEQ!�*�*�@�OS��l4� 4�60ENABy� PTION�3��r���^GCF�!� �@60J�Q���R�d!��G�P�EDIT�� ��� ��KAQ"� �E�(�NU'(AUT<Y�%COPYAQ�(2,�qe�M�N< @+^��PRUTm� C"�N�OU�2$G���$��RGADJZ��u2X_��IX�P���&���&W�(P�(�~��&9�� 
�N�P_�CYCy�v�RG�NSc�{�s�LG�O£�NYQ_FREQSrW@��X1�4�L�@�2P0�!�c@�"�CRE��Mà�IF�q�NA���%�4_Gf�STA�TU~�f��MAI�L��|CIq�=LA�ST�1a*4ELE�Mg� ��QrFEASIt;�ւΰ ��B"�F�AF����I� ��O2�E u�&vBAB��PE� =��VA�FzQ�I��TqU�[��R��S�FRMS_TRpC�Qc���C��Z�
��1�D �Ens؆�	MB 2� `���N� 3V�R2WR*���шR8^W�wj�DOU�^��N�,2PR`�hٞ1GRID��B7ARS!�TYu�r�Op�� |E_�4!� �R�TO��>d� � �����POR�c~vbS�RV�0)"dfDI[�T�`;aNd�pXg
��Xg4Vi��Xg6Vi7�Vi8:aZFʒg�~z $VALU�C�0�3D1@v�F05��� !pT���S�1-ȆAN/��b�1�R�]11ATOTA�L����=sPWE3I|�QStREGENQzfr��X�H�]5	v�( TR�CS�Qq_S3��wfp�V�!��r��BE�3�PG0B��( sV_H�PDA8(��p�S_Ya����i6S��AR(�2�� �"IG_SE��3�pb�5_� �tC=_�V$CMPl��KDEp�G���Iš�Z~�X��R�aENH�ANC.� p� Qr�2���IN�T9`cq�F���M�ASK�3�@OVRMP �PD�1-��W�aХT�l�_RF|�{�V�PSLGP�
g�9�j5��,��;pDpS���4��aU���n �TE����`���`k���Jx^�Y�y3IL_Mx40�s��p��TQ( �P��@����V.�C<��P_ �R�F�M]�V�1\�V1j�2y�2�j�3y�3j�4y�4 j���p۲������vܲIN�VIB8�P6�#��*�2&�22�U3&�32�4&�42���6�|�J�  �T $MC_FK `� �L>�J�х�1pMj�Iу��zS ���1���KEEP_HNADD���!鴓@�C��0 	��Q����
�O!��v ���p
�և
�REM!�	�Cq�RF�]��b�U�4e	�HPW�D  �SB�M���PCOLLAAB*�p��/q�2cIT/0��Q"NO1�FCALp⎵��� , �FLv�AO$SYN���M���Ck��RpUP_D�LY��zDEL�A9�Dq�2Y AD�(��aQSKIPNO�� �`� O��cNT����c�P_�  ��׾ ��cp���q�� ���o`��|`�ډ`��@�`�ڣ`�ڰ`��9�!O�J2R0  �lX�@TR3H��1AH��� �H���v�RD�Cq��� � R"�R, 5��R�1��8E��5TRGE�_C��RFLG"���9W�5TSPC�1�UM_H��2TH�2N}Q�;� ?1� ��;��Q>02 � D� ˈ<��@2_PC3W��S���1Y0L10_�Cw2 ,��� � $\� U@�� V7�����0��VU\����� rd���C6�,��7��DrZ Gs�RUVL1[��1h���10]�_�DS����ʑ�PK 11�� lڰ����q��AT?��$�Q [7�R��K 5T����HOME� _2h�n������&0`3h����!3E ��c4h�hz����� �`5h���	//-/?/W `6h�b/@t/�/�/�/�/�'7h��/�/??'?9?W8h�\?n?�?�?�?v�? *�FPS��>��  �Aa�{p���_�Ed�� T=�nD4vnCIO�䑎II@`�O��_�OP�E�C.r��]P�OWE	�� �X@�f�	�$�$Cd�S����i��A3�3� �@��SI��G�P0�QIRT�UAL�O
QAAV�M_WRK 2 �7U 0  �5Q�n_zXk_�] ��\	[ �]�_3�8P��_�_�Ve�\#m/o��Q5ojo|o�dHPBS��� 1Y� <Xo�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯�ݯ�bC$�AXLM��@���c  �d�IN����P+RE
�E�J�-�'_UP��[�7QHP?IOCNV_��k �	�Pr�US>��g�cIO)�V 1]U[P $E`��Q0ս9lҿ8P?�� � ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o�o�o�o�m�LAR�MRECOV �a��-���LMD/G ��ɰ��LM_IF  ���ை����z�v���%�6�, 
 6�_��r� ��������̍$w��� ׏��8�J�\�n�����NGTOL  �a� 	 A �  ��ț�PPI�NFO ={� <v����1��  I�3�a�"rP��� t��������ί���>�o����j�|��� ����Ŀֿ������0�B�PzPPLIC�ATION ?����+��HandlingTool ��� 
V9.30�P/04ǐM�
�88340�å�F90����202�ť�|�Ϭ�7DF3���M̎�NoneM��FRAM� �6��Z�_ACTI�VE�b  sï� � p�UTOMO�Dz�A���m�CH�GAPONL�� ���OUPLEDw 1ey� �������g�CURE�Q 1	e{  T*���	p��xw���#r�g���e�HN����{�HTTHK)Y��$r��\[�m� ���O�	�'�-�?�Q� c�u����������� ��#);M_q ������ %7I[m� ��/���/!/ 3/E/W/i/{/�/�/�/ ?�/�/�/??/?A? S?e?w?�?�?�?O�? �?�?OO+O=OOOaO sO�O�O�O_�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q��c���1�TO��|��p�DO_CLEA�N��n��NM  �� �B�T��f�x���%�DSPDgRYR��m�HI���@/�����,�>� P�b�t���������ίj�MAXa�ۄ�������Xۄ������p�PLUGG��܇�Ӯ��PRC��B�" ��ׯF�OK���^ȔSEGF��K�� �����.�����,�8>�v���LAPӟ� ��Ϥ϶��������π�"�4�F�X�j߯�T�OTAL�7���U�SENUӰ�� ����ߖ�1�RGDI_SPMMC����C����@@Ȓ��O�ѐ�����_STRING 1
�ۿ
�M��S�l�
A�_ITE;M1K�  nl�g� y������������ 	��-�?�Q�c�u����������I/O SIGNALE��Tryout� ModeL�I�np��Simul�atedP�Ou�tOVER�RА = 100�O�In cyc�lP�Prog� AborP�~��StatusN��	Heartbe�atJ�MH F�aul��Aler�	�������*<N`  ׃G�ׁY�c��� ��////A/S/e/ w/�/�/�/�/�/�/�/wWOR��G�-1� ?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO�cOuO�O�O�NPO E��@E;�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8oJo�BDEV�Nu`�O bo�o�o�o�o�o�o ,>Pbt�������PALT��E?�A�S� e�w���������я� ����+�=�O�a�s����GRI�G뽑 1������	��-�?� Q�c�u���������ϯ�����)�����R �a�՟;��������� ѿ�����+�=�O� a�sυϗϩϻ���O�PREG��y��� -�?�Q�c�u߇ߙ߫� ����������)�;��M�_�q����$AR�G_-0D ?	��������  	$���	[��]���������SBN_CONFIG���� ��CII�_SAVE  ���)���TCEL�LSETUP ���%  OME�_IO����%M�OV_Hn�����R�EPd�����UTO/BACKY���#�FRA:\��� ����)�'`rl ��&� 7�"� 24�/06{  09:_35:24������͓����� �+=Oas��������� �/1/C/U/g/y/�/ /�/�/�/�/�/	?�/ -???Q?c?u?�?�?p�ׁ  _��_\�ATBCKCTL.TM���?�?�?O\ O��INI�Y��-���MESSA�G9�GA)��RKODGE_Ds�<��zH�Ow`�O��PAUS��@ !��� ,,		�����O �G�O__#_%_7_q_ [_�__�_�_�_�_�_��_%o���D�@TSK  �M&,O���UPDT�@EGd��`�FXWZD_E�NBED��fSTApDE��e��XIS�?UNT 2��&��(�� 	 �6G0 �8/� 0�=�y� �����Tpp�p�p�p��GA7qUg~)qq��~�ĥS�,��[ �?t� {!jD�ph���fMETc��2LfE� P q@��n�A1�A��"A�A�$)BhS�}�=���>�g��>�F?O`��>�k^>�����}SCRDCFG� 1�� �A�&������@ԏ�����Q=� ��H�Z�l�~�����	� Ɵ-����� �2�D�0��域���GR�`�`X�O���0NA����s	��_EDC@�1n�� 
 ��%-�0EDT- q����%�,q�I�(��������������  ����2����*���bB���@*�q���ϧ���3b� ��@Ͻϯd?�����=�O���sϏ�4.ߞ�{� ����W���	�߱�?���5��j�G����#�@������}�6�� 6��Z�����Z����I��7�����&� �λ�&m������!8^ҿ����	͇@�9K�o��9*�w��	�S�0�;��CR���� B/T//�/��w/�/��РNO_DE�L����GE_UN�USE���IGALLOW 1���   (*SYSTEM*�s�	$SERV_�GR�;B0�@REG�K5$m3�|B0NU�Mp:�3�=PMU|� �uLAY�p��|PMPA�LD@�5CYC10��.�>�0�>CUL�SU�?�=�2�AM3�LOWDBOXOR=It5CUR_D@�=�PMCNV�6�D@10�>�@T4�DLI�`=O_9	*�PROGRAJ4?PG_MI�>�OFPAL�E_UP�B7_B>$FLU?I_RESU�7p_z?�_�TMRY>1p�,�/�b�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv����������"LAL_OUT 1;l���WD_ABOR�0�?d�ITR_RT/N  �����g�?NONSTOǠ��� 8CE_RIgA_I0��ۀ���ŀFCFG ���۔���_L�IMY22ګ �  � 	i�DJ��<e�g��5��P� 9���������a
���u��PAQP�GP 1������Q�c�u�4�CXK0����C1��9��i@���PC��CV��U]��d��l��s��XP���C[٤m���v���������W C����-�����?�ÂHE� ON�FI�Pq�G�G_Pv�@1� �% �������ǿٿ���|�G�KPAUSaA31�ۃ �B� W��Eσ�iϓϹϟ� ���������#�I�/ߠm��eߣ��M��N�FO 1"��� �7��ߖ���B��L���A��=AV�������� ¶��C��y�C�K���3�����B����4�F�ŀO��c�COLL/ECT_�"�[�����EN�@��y���nk�NDE��"��3�"1234?567890�� \1�� ��֕H&��)M�r�\,L�^���]+ ������������C  2�Vhz�� ����
c. @R�v����t����� ��>��IO !���q���u/�/�/�/C'[TR�2"'-(�Pb^)
��.R�#R-x�*W� 9_MOR�$� �;�l5��l9 �?r?�?�?�?�;E2�*�%S=,W�?@�@�I�C�PK)DցC��R�&u�XOWAWBC_4  A�q���P�x�PA"@Cz + B�@CG�B8��A�C  @yB���Pց:d�43? <#�
�E��P�I�O�C=AI��'GM�?�C�(S=���Qd�=AT_DEFPR/OG �;%�/m_|APINUSE��V�ۅ�TKEY_TOBL  s�ہ����	
�� �!"#$%&'()*+,-./��:;<=>?@A�BCDPGHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������Ga���͓���������������������������������耇���������������������$��PLCK�\���P΋PSTAn��T_A�UTO_DO��NFsIND���n���R_T1wT2�N����5ŀTRL^CPLETE���z�_SCREEN ��kcs�cÂU��MMEN�U 1)O� < �[_#�q��,�a��� >�d���t���ӏ���� 	�����Q�(�:��� ^�p�������̟�ܟ �;��$�q�H�Z��� �������Ưد%��� �4�m�D�V���z��� ٿ��¿�!���
�W� .�@ύ�d�vϜ��Ϭ� �������A��*�P� ��`�r߿ߖߨ����� ���=��&�s�J�\� �����������'��,�p_MANUAL�EqDB
12�v��iDBG_ERR�LIP*�{h! �0�������g�N_UMLIM�s:Q�OE�@DBPXWO_RK 1+�{���>Pbt��-DBwTB_�q ,���kC3!VD!DB__AWAYo�h!oGCP OB=��A�_AL���o�k�Y�p�uO@`�_�� +1-�+@
-k�-6[��_M+pI�S�`�@"@�ON�TIM�w�ODɼ�&
�U;MO�TNEND�_:R�ECORD 13��{ ��[CG�O�f!T/[K��/�/ �/�/_(�/�/f/?�/ ??Q?c?�/?�??�? ,?�?�?OO�?;O�? _O�?�O�O�O�O(O�O LO_pO%_7_I_[_�O _�O�__�_�_�_�_ l_!o�_,o�_io{o�o �oo�o2o�oVo /A�oeP^�
 ���R���=� �a�s��������*� ߏN���'���ԏ]� ̏��������ɟ۟v� ��n�#���G�Y�k�}����TOLERE�NC�B�0� L���g�CSS_C�NSTCY 24J	�t���.�� ����0�>�P�b�x� ��������ο�����(�:�äDEVI�CE 25ӫ ��ϟϱ������π����/�AߟģHNDGD 6ӫ�� CzT�.!ơLS 27t�S����߀������/�U�ŢPARAM 8G�b�A�Ք�RBTw 2:8��<���CkA�� ·�  �� A���.S�B���A�B�  ���������.�� ����A�A�C����c�u�l���C�A�D�(�k�pz�A�A��HA�c��A�	�? (uL^p��|�A�Bt/�D���C��_ 	 �A=��ABffA#33AҊ���A�A�C%f��a��A�J���7B]��B��BffBᴠ�33C$.@R� ( ���A� ����
/��// )/;/�/_/q/�/�/�/ �/�/�/�/<??%?r? I?[?m??�?�?�?�? �?&O8O�PObOMO�O qO�O�O�O�O�O_� OOL_#_5_�_Y_k_ �_�_�_�_ o�_�_6o ooloCoUogo�o�o �o�o�o�o �o	 h�O�w���� �
��.�	__I'� 1_�q��������ˏ ݏ���%�r�I�[� ���������ǟٟ&� ���\�3�E�W���� ȯ���ׯ�"��F� 1�j�E�s�����m��� ����ѿ�0���f� =�O�a�sυϗ��ϻ� �������'�9�K� ��o߁�����[���� (��L�7�p��m�� ������������$��� ��l�C�U���y��� �������� ��	V -?�cu��� �
��@+dO �s������� �*///`/7/I/[/ m//�/�/�/�/?�/ �/?!?3?E?�?i?{? �?�?�?�?�?�?�?FO �jOUOgO�O�O�O�O �O�O__�'O9OO =_O_�_s_�_�_�_�_ �_�_�_oPo'o9o�o ]ooo�o�o�o�o�o �o:#5��O� ���� ��$���H�Fz�$DCSS�_SLAVE �;���w���`�_4D � w���AR_M�ENU <w�  >�؏���� �2�^r�Ǐ\�n�\���SH�OW 2=w� � fr[q����Ə �����,�>�D�b�t��� ����ҟϯ� ���)�P�M�_�q� ��������˿ݿ�� �:�7�I�[ς�|Ϧ� �ϵ���������$�!� 3�E�l�fߐύߟ߱� ���������/�V� P�z�w������� ������@�:�d�a� s�����������\��� *�H�N�K]o� �������2 8�GYk}�� ����"�1/ C/U/g/y/�/��/�/ �/��//?-???Q? c?u?�/�?�?�?�/�? ?OO)O;OMO_O�? �O�O�O�?�O�?�O_ _%_7_I_pOm__�_ �O�_�O�_�_�_o!o 3oZ_Woio{o�_�o�_ �o�o�o�oDo- Se�o��o��� ���.�=�O����CFG >������q��dM�C:\��L%04�d.CSV\��pc��������A ՃCH݀z�v�w�#�
�q���:�J�8�<7���JP�j�)��́�p+�n�RC_OUT ?z������a�_C_FSI ?��? |�� ���@�;�M�_��� ������Я˯ݯ�� �%�7�`�[�m���� ����ǿ�����8� 3�E�Wπ�{ύϟ��� ���������/�X� S�e�wߠߛ߭߿��� �����0�+�=�O�x� s����������� ��'�P�K�]�o��� ��������������( #5Gpk}�� ��� �H CUg����� ��� //-/?/h/ c/u/�/�/�/�/�/�/ �/??@?;?M?_?�? �?�?�?�?�?�?�?O O%O7O`O[OmOO�O �O�O�O�O�O�O_8_ 3_E_W_�_{_�_�_�_ �_�_�_ooo/oXo Soeowo�o�o�o�o�o �o�o0+=Ox s������� ��'�P�K�]�o��� ��������ۏ���(� #�5�G�p�k�}����� ��şן �����H� C�U�g���������د ӯ��� ��-�?�h� c�u���������Ͽ�� ���@�;�M�_ψ� �ϕϧ���������� �%�7�`�[�m�ߨ� �ߵ����������8� 3�E�W��{����� ���������/�X� S�e�w����������� ����0+=Ox s������ 'PK]o� �������(/ #/5/G/p/k/}/�/�/ �/�/�/ ?�/??H?�C?U3�$DCS_�C_FSO ?�����1? P [?U? �?�?�?�?�?O
OO .OWOROdOvO�O�O�O �O�O�O�O_/_*_<_ N_w_r_�_�_�_�_�_ �_ooo&oOoJo\o no�o�o�o�o�o�o�o �o'"4Foj| �������� �G�B�T�f������� ��׏ҏ�����,� >�g�b�t��������� Ο�����?�:�L� ^���������ϯʯܯ�g?C_RPI~> �?�;�d�_�
�}?.�`p����ݿj>SL�@���9�b�]�oρ� �ϥϷ���������� :�5�G�Y߂�}ߏߡ� �����������1� Z�U�g�y������ ������	�2�-�?�Q� z�u������������� 
)RM_q ������� *%7Irm� ����/�ϛ� ,�/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO sO�O�O�O�O�O�O_ __'_P_K_]_o_�_ �_�_�_�_�_�_�_(o #o5oGopoko}o�o�o �o�o�o �oH CUg��������� ����NOCODE @������PR�E_CHK B쟻3�A 3��< �7�����<���� 	 <��� ��?#ۏ%�7��[�m� G�Y�������ٟ�ş �!����W�i�C��� ��y�ïկˏ���� ��A�S�-�_���c�u� ��ѿ�������=� �)�sυ�_ϩϻϕ� �������'�9���E� o�I�[ߥ߷ߑ����� ����#����Y�k�E� ���{�������� ���C�U��=����� w���������	���� ?Q+u�a�� ����); _qg�Y��S� ���%/�/[/m/ G/�/�/}/�/�/�/�/ ?!?�/E?W?1?c?�? ���?�?o?�?O�? �?AOSO-OwO�OcO�O �O�O�O�O_�O+_=_ _I_s_M___�_�_�_ �_�_�?�_'o9oo]o ooIo�o�oo�o�o�o �o#�oGY3E ��{����� o�C�U��y���e� ����������	��-� ?��K�u�O�a����� ����͟��)��1� _�q��}�������ݯ �ɯ�%���1�[�5� G�����}�ǿٿ��� ����E�W�1�{ύ� G�u����ϯ������ /�A��-�w߉�c߭� �ߙ���������+�=� �a�s�M���ϑ� ������'��3�]� 7�I������������ ������GY3} �i������� �C/y�e �������-/ ?//c/u/O/�/�/�/ �/�/�/�/?)?�? _?q?K?�?�?�?�?�? �?�?O%O�?IO[O5O O�OkO}O�O�O�O�O _�O3_E_;?-_{_�_ '_�_�_�_�_�_�_�_ /oAooeowoQo�o�o �o�o�o�o�o+ 7aW_i_��C� ����'��K�]� 7�i���m��ɏۏ�� �����G�!�3�}� ��i���ş����� �1�C��g�y�S�e� ���������ѯ�-� ��c�u�O������� Ͽ�ןɿ�)�ÿM� _�9�kϕ�oρ����� �������I�#�5� ߑ�kߵ��ߡ����� ��3�E���Q�{�U� g������������ /�	��e�w�Q����� ����������+ Oa�I���� ���K] 7��m���� �/�5/G/!/k/}/ se/�/�/_/�/�/�/ ?1???g?y?S?�? �?�?�?�?�?�?O-O OQOcO=OoO�O�/�/ �O�O{O�O_�O_M_ __9_�_�_o_�_�_�_ �_oo�_7oIo#oUo oYoko�o�o�o�o�o �O�o3Ei{U �������� /�	�S�e�?�Q����� ��я㏽���� O�a�������q���͟ �������9�K�%� W���[�m���ɯ��� ��ٯ�5�+�=�k�}� ������������տ �1��=�g�A�Sϝ� �ω����Ͽ��������Q�c����$D�CS_SGN �CS�����g��06-JU�N-24 12:�37 EӘ�09:�39������ _X�L���������������#M���M��Þ�ǧj�����{�VE�RSION ���V4.2.�10�EFLOG�IC 1DS���  	�D���X�k�X�z�M�P�ROG_ENB � ��b��Л�U?LSE  ����M�_ACCLI�M��������WRSTJNT�����w�EMO���ѷ�L��INIOT EZ�O���OPT_SL ?�	S�1�
 	�R575�Ӆ�74*��6��7��5A��1��2��l���G�h�TO  t���.�H�V?�DEX��d����FPATHw A��A\4����HCP_CLNTID ?+�b� l������IAG_GRP� 2JS�� �a[��D�  D�� �D  B�  ;B�@ff��/CB�@[��W�@��q��B�N��C�-Bz�w�Bp@e`���mp3m7 �78901234�56�*�[�� � Ao�mAj�1AdA]��
AW|�AP��AJ-AC�/A;�A4�H���@�  Aʩ�A�A3!_A�@@��B4��� ��t���
�u�ƨApffAj��yAeK�A_��AY��AS�� MC�AF��A@ �O�+/=/O$�O�c K�w(@�X�?8��@��y�/�/�/�/�/8��;d�2�5?@~�ff@x1'@q���@kC�@d��D@]��@Vv�6?H?Z?l?~?8�s�0l��@e���@^��@W\)@O��@H�0�?<@7K�@.V��?�?�?�?
O8S�@M00G<@A���@<1@5���@/l�@(�Ĝ@!�0�\ NO`OrO�O�Ox'g�L_ K�;_�_�__g_�_�_ �_�_o�_�_�_Yoko@Io�o�o+o�oX�"�� 2�17A�@J>���R
q?�33?wY��r��J�7'Ŭ2q63p4w�F>r��LJ�@�p�Zr�
=�@�@�Q�jq��@G Ah�@���@�T= c<���]>*�H>�V>�3�>����J<���C<�p�q�x��� ��?� �C� � <(�U�� 4Vr�33��@
���A@��?R�oD� �mR�x���Q��t�����Z�Џ��؏�,��i?��7N�>�(�y>�@Z�=���Jo��G�v�G�J �B�E�����a��@ǐ�@���@��@OQ�?L ���ŲI�P���&�
��'��@�K�����Ag�q�PC�  ?C���Cuy�
����ʯ ?մ�}Q�?S̑?ˤ�?)5�
����m��Ľ��¶�MC�x_�C�L8��>(����4���X��v����*
��3������F�ǿB���ֿ����E�t�9���þ��<>K`.>�?YؾHܹ
�I����CT_CON�FIG K|3���eg���STBF_TTS��
����"�����:��{�MAU��~�MSW_CF���L  K �OCoVIEW	�MI�U����߭߿��� �������0�B�T� f�x���������� ����,�>�P�b�t� ������������� ��(:L^p� ����� � 6HZl~�������/��RCB�N��!�X.F/ {/j/�/�/�/�/�/���SBL_FAUL�T O9*^�1G�PMSK��7��TDIAG P���Uѵ����q�UD1: 6789012345q2�q���%P�ϭ?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O ��a6�I'�
�?_��TORECPJ?\:
j4 \_�7u[�?�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�O�O_� _�UMP_OP�TION��>qT�RB���9;uPM�E��.Y_TEM�P  È�33B����p�A�pyt�UNI'��ŏq6�Y�N_BRK Q�t�_�EDITOR� q&qh�r_2PEN�T 1R9) � ,&MAIN� BARRA_E?STEIRA����&PEGA_%��b�&COLO�CO��pNO^����&PICK1_PLACE0 ���?���P�PRENS�]��&SUM#IR~��D�Ѓ����?���UP~�@�&T�W���s��/��������Ο��� A�(�e�L��������� �����ܯ� �=�$��6�s�Z��pMGDI_STA�u~��q�u�NC_INFO �1SI��b��������Կⷮ���1TI� ��o#��G�
G�d�o}Ϗϡϳ� ����������1�C� U�g�yߋߝ߯����� ����Hu� �2�D�R� j�R�x�������� ������,�>�P�b� t�������������Z� �#5Ga�k} ������� 1CUgy�� ������	//-/ ?/Yc/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? ��?O%O7OQ/GOmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�?Ooo /o�_[Oeowo�o�o�o �o�o�o�o+= Oas����� �_�_��'�9�So]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�K�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�C�5� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ�������� �!�;�M�W�i�{�� ������������� /�A�S�e�w������� ��������+E� Oas����� ��'9K] o����1��� �/#/=G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?��?�?	OO5/ ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�?�_ �_oo-O#oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���_�_���� 7oA�S�e�w������� ��я�����+�=� O�a�s��������� ߟ���/�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������͟׿���� '�1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߫�ſ ���������;�M� _�q��������� ����%�7�I�[�m� ������߯������� �)�3EWi{� ������ /ASew���� �����/!+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?/��?�?�? �?/#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �?�_�_�_�_Oo-o ?oQocouo�o�o�o�o �o�o�o);M _q���_��� �	o�%�7�I�[�m� �������Ǐُ��� �!�3�E�W�i�{��� ��ß՟矝��� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}� �ߩ����������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u����߫��� ��������);M _q������ �%7I[m �������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?���? �?�?�?�OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�?�?�_�_�_�_�? �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�_� ����_�	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q��y�����˟� ۟��%�7�I�[�m� �������ǯٯ�����!�3�E�W�i��� ��$ENETMO�DE 1U��  ���������»��R�ROR_PROG %��%������TABLE  ���Q�c�uσ���SEV_NUM� ��  �������_AUT�O_ENB  �̵��ݴ_NO�� �V������ W *���������	�����+���(�:ߞ��FLTR����H�IS�Ð�����_A�LM 1W�� e����̍�+;߀��������0�?�_\����  �����²u꒰TCP_V_ER !��!���@�$EXTLOGo_REQv�������SIZ����ST�K�������T�OL  ��Dz�~��A ��_BWDU�*�Z�V�ǲ?�DID� X��Z�����[�ST�EPl�~�����OP�_DO���FAC�TORY_TUN�v�d��DR_GR�P 1Y��`�d �	p�.° �*�u���RH�B ��2 ���� �e9 ����bt� A���aA�c�B���pBy.A��HGBn�@���-AS�*B�@:�A+A�^�B]�� ���
C.g�R  A]M@��W�@L�f?�v��u
 IǍo����@���u��a[ /��$/�B�  F!Aݠ��33R"�3]3�UUTn*@�� /ȷ>u.�>*��<��Ǌ�E�� F@ ξ"�5W�%�J���NJk�I'�PKHu��IP��sF!���?�  ?�/9��<9�8�96C'6<�,5������1|�+��E�� � f�e��M��F�EATURE �Z�V�Ʊ�Handling�Tool �5���English� Diction�ary�74D S�t�0ard�6�5A�nalog I/�O�7�7gle S�hift Outo� Softwar�e Update�%Imatic B�ackup�9SAg�round Ed�it�0�7Came�ra�0F�?Cnr�RndImXC�Lo�mmon cal�ib UI�C�Fn�qA�@Monito�r�Ktr�0Rel�iab@�8DHC�P�IZata A�cquis�CYiagnosOA�1[�ocument �Viewe�BWu�al Check Safety�A~�6hanced�F4�:�UsnPFr�@�7�xt. DIO ��@fiRT�Wend.�PErr�@LQR�]J�Ws�Yr�0�P E���:FCTN Me�nu�Pv S8gTPw In'`facNe�5GigE`nrej@�p Mask Ekxc�Pg�WHT^`�Proxy Sv�oT�figh-Spe�PSki�D�eJP~�PmmunicN@7ons�hurE`'`�_�1abconne�ct 2xncr``stru�2z>p�eeQPJQU�4KA�REL Cmd.� L�`ua�husR�un-Ti�PEnyvkx(`el +R@�sP@S/W�7License�Sn\�P�Book(Sys�tem)�:MAC�ROs,�b/Of'fse@�uH�P8@�_�pMR�@�BP^MechStop�at.p6R�ui�RKj�ax�P�0P@)�od@witch��>�EQy.���OptmЏ�>��`filn\=�g�w�uulti-T��`tC�9PCM funHwF�o3T�R?�^f�Regi�pr�`I�rigPFV����0Num Selb�|���P Adju�`��J�tatu�
�iZ�5RDM �Robot�0scgove�1F�ea7���PFreq An;ly�gRem`��Q�n�7F�R�Serv�o�P���8SNPX� b�rNSN^`C�lifQɮBLibr�3鯢0 q������o�ptE`ssag?��4�� -C��;���/I_mB�MILI�Bk�E�P Fir�m6BU�PEcAcc<k@sKTPTX_C�eln���F��1��V�orqu@imGula�A�A�u���Pa�qU�j@�Ã&ε`ev.B�.@ri�P޿USB poort �@iP�P�agP��R EVN�T�ϗ�nexcept�P��t��ſX�]�VC�Ar�b�bf�V@2PҦ�$����SܠsSCصV�SGEk��a�UI�;Web Pl!��ާ��Խ`��TeQfZDT Appl�d�:�ƺ� ��GridV�pla�y�R�WD4�R
�.��:n�EQ+��r-10�iA/7L*��1G?raphic���5�dv�SDCSJ�c�k�q�5larm �Cause/��e}d�8Ascii�a���LoadnP�U�pl,�Ol�0�AG�u�6N�`���yFyc�@�r�����PV��Jo��m� c�R���c���m�./�����Q�2*u:eRAJ��P�ٌ�4eqinL����8N�RT��9On�0e Hel�HJ�`oI�alletiz?��H�����_�tr�[R?OS Eth�q���T@e�ׅ�!�n�%�2D�tPkg&�Upg~�(2D�V-�3D Tr�i-jQEAưDe�f.qEBa)pde`i��� �bImπqF�f��nsp.q�=�464MB D�RAMZ,#FRO�5/@ell�<�Mshf!r/�'c%3@YpLƖ,ty@s˒xG��m��.[�� ���BU���Q�B�=mai�P߫�]Q����@q6wlu����^`�x�R�?eL� Sup�������0�P�`cr ��@�R���b䚮�pr1ouest�rt~QQ��ߋL!�4O��q�$�K��l Bu�i7�n��APLCdOO�EVl%��CGUN�OCRG�O��DR���O
TLS_��BU�/_��K�qN_d�TA�OxVB�_�W�ܑZ���_TCB�_�V�_�W���WF+o�V�O�W._8�W�ņoTEH�o�f0�O�gt�oTEj�xV!F�_w�_xVGoTw�BTw~oxVH�xVIaA��v�xVLN�yUMz�bo�f_xV	N�xVP���^xV	R&xVS��܇ʏ���W��v���VGF:�L�P2_h��h��V�h��_g�D��h�F0Foh��g�RD�� 7TUT��01:�L�y2V�L�TBGG���v�rain�UI���
%HMI���p#on��m�f�"��F�&KAREL9� �TPj��<6� SWIMEST&ڢF0O�<5�
"a� X�j�������ͿĿֿ ���'��0�]�T�f� �ϊϜ����������� #��,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ ����������$�Q� H�Z���~��������� ���� MDV �z������ 
I@Rv ������// /E/</N/{/r/�/�/ �/�/�/�/???A? 8?J?w?n?�?�?�?�? �?�?O�?O=O4OFO sOjO|O�O�O�O�O�O _�O_9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l���������Ə ����)� �2�_�V� h����������� ��%��.�[�R�d��� ������������!� �*�W�N�`������� �����޿���&� S�J�\ωπϒϤ϶� ��������"�O�F� X߅�|ߎߠ߲����� �����K�B�T�� x����������� ��G�>�P�}�t��� ���������� C:Lyp��� ���	 ?6 Hul~���� �/�/;/2/D/q/ h/z/�/�/�/�/�/? �/
?7?.?@?m?d?v? �?�?�?�?�?�?�?O 3O*O<OiO`OrO�O�O �O�O�O�O�O_/_&_ 8_e_\_n_�_�_�_�_ �_�_�_�_+o"o4oao Xojo|o�o�o�o�o�o �o�o'0]Tf x������� #��,�Y�P�b�t��� ������������ (�U�L�^�p������� ���ܟ���$�Q� H�Z�l�~�������� د��� �M�D�V��h���  �H552}���21n��R78��50���J614��ATU]PͶ545͸6���VCAM��CRIn�UIFͷ28	ƷNRE��52��R�63��SCH��DwOCV]�CSU���869ͷ0ضEI�OC9�4��R69���ESET���J�7��R68��MA{SK��PRXY!�]7��OCO��3�h����̸3�J6˸�53��H2�LCH^��OPLG�0֯MHCR��S{�MkCS�0��55ض�MDSW���OP��MPR�M�@�0n̶PCM �R0���ض��@�51�5u1<�0�PRS�ǻ69�FRD�FwREQ��MCN��{93̶SNBAE�^3�SHLB��M��tM���2̶HTC��TMIL����TP�A��TPTX��EL��Ѐ�8������wJ95,�TUT׻95�UEV��U�EC��UFR�V�CC��O��VIP��CSC,�CSGt8�r�I��WEB�7HTT�R6C�N��CGIG��IP�GS)RC�DG��H77��6ضR�85��R66�Ru7��R:�R530�K680�2�q�J��*H�6<�6,�RJح�j0�4�6o64\��5�NVD��R6��R84Tg�����8�90\���J9&3�91� 7+����,�D0oF�CL9I���CMS�� n�STY��TO䶴q���7�NN�O�RS��J% ��j�O]L(END��L���Sf(FVR��V3�D���PBV,�A�PL��APV�C�CG�CCR|�C�D��CDL@CS�Bt�CSK��CT�CTBL9��U0,(�C��y0L8C��TC� �y0�'TC(7TC���CTE\��07T�Eh��0��TFd8FJ,(GL8GI�8H�8�I��E@�87�CTM�,(M�8M@8N�8P�HHPL8Rd8(TSrd8W�I@VGF�GP2��P2���@�H�{7VPD�HF �V�PSGVPR�&VT���YP��VTB7Vs�IH��VI aH'�VK��VGene�����_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 I[m���� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/?�?+?=?O?a?s?�?�  H55�hT�1�1[U�3R78��<50�9J614έ9ATU�T�454u5�<6�9VCA�Dn�3CRI,KUI8Tv�528-JNRE�:�52JR63�;S{CH�9DOCV�J�CU�4869�;0N�:EIO�TsE4�:�R69JESET��;KJ7KR68ތJMASK�9PR�XYML7�:OCOB\3�<�J)P�<3|Z[J6�<53�JH�\�LCH\ZOPLGz�;0�ZMHCR]Z]SkMCS�<0,[{55�:MDSW}kv�[OP�[MPR�Zt�@�\0�:PCMLJ�R0�k)P�:)`�[5�1K51|0JP�RS[69|ZFR�D<JFREQ�:M�CN�:93�:SN�BA}K�[SHLB��zM�{�@ll2�:H{TC�:TMIL�<��JTPA�JTPT�X�EL�z)`�K8��;�0�JJ95\JT�UT�[95|ZUE�VZUEC\ZUF]R<JVCC��O<jwVIP,�CSC\��CSGlJ�@I�9W�EB�:HTT�:R�6{L��CG{�IG�[�IPGS��RCv,�DG�[H77�<�6�:R85�JR6�6JR7[R|R[53{68|2�ZR�@Jml,|6|6\JQR�\	P|4L�6��64��5�kNVDvZR6+kR84<�h��IP,�8��90��6�KJ9�\91��̫�7[KIP\JD0�F���CLI�lKCMqS�J9��:STY,��TO�:�@�K7�LN]N|ZORS<jJ���MZZ|OLK�END�:L�S��FVR��JV3D,�KKPB�V\�APL�JAP�V�ZCCG�:CC�RjCD�CDL�̚CSB�JCSKv�jCTK�CTB�݈\���\�C�z���C�L�TCLJ�l�TCv��TCZCTE�J���|�TE�J��<�TUF��F\�G��G��
l�Hl�I�z)�l�k�WCTM\�M\�M��UNl�P,�P��R�ܖ;�TS��W��̚V�GF��P2��P2p�z �VPD�FLJVP;�VPR���VT�;� �JVT�B��V�KIH�VXِM�<�VK,�V{�Gene�8�83E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ��������� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ��������1�C�U� g�y������������� ��	-?Qcu ������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ �/�/�/�/?!?3?E?�W?i?{?�7�0�STD�4LANG�4�9�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~��������� �2�D�V�RB=T�6OPTNm�� ������Ǐُ���� !�3�E�W�i�{�����8��ß�5DPN�4� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G��Y�k�}ߏߡ߳�ted �4�8������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u��������� ������);M _q������ �%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ������*�<�N�`�r�99���$F�EAT_ADD �?	�����~��  	�� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu������DEMO �Z��   ���}��'��0� ]�T�f����������� ����#��,�Y�P� b�������������� ���(�U�L�^��� ���������ܯ�� �$�Q�H�Z���~��� �����ؿ��� � M�D�Vσ�zόϦϰ� �������
��I�@� R��v߈ߢ߬����� �����E�<�N�{� r����������� ��A�8�J�w�n��� ������������ =4Fsj|�� ����90 Bofx���� ���/5/,/>/k/ b/t/�/�/�/�/�/�/ �/?1?(?:?g?^?p? �?�?�?�?�?�?�? O -O$O6OcOZOlO�O�O �O�O�O�O�O�O)_ _ 2___V_h_�_�_�_�_ �_�_�_�_%oo.o[o Rodo~o�o�o�o�o�o �o�o!*WN` z������� ��&�S�J�\�v��� �������ڏ��� "�O�F�X�r�|����� ��ߟ֟����K� B�T�n�x�������ۯ ү����G�>�P� j�t�������׿ο� ���C�:�L�f�p� �ϔϦ�������	� � �?�6�H�b�lߙߐ� ������������;� 2�D�^�h������ �������
�7�.�@� Z�d������������� ����3*<V` �������� /&8R\�� �������+/ "/4/N/X/�/|/�/�/ �/�/�/�/�/'??0? J?T?�?x?�?�?�?�? �?�?�?#OO,OFOPO }OtO�O�O�O�O�O�O �O__(_B_L_y_p_ �_�_�_�_�_�_�_o o$o>oHouolo~o�o �o�o�o�o�o  :Dqhz��� ����
��6�@� m�d�v�������ُЏ ����2�<�i�`� r�������՟̟ޟ� ��.�8�e�\�n��� ����ѯȯگ���� *�4�a�X�j������� ͿĿֿ����&�0� ]�T�fϓϊϜ����� �������"�,�Y�P� bߏ߆ߘ��߼����� ����(�U�L�^�� ������������ � �$�Q�H�Z���~��� ������������  MDV�z��� ����I@ Rv����� ��//E/</N/{/ r/�/�/�/�/�/�/�/ 
??A?8?J?w?n?�? �?�?�?�?�?�?OO =O4OFOsOjO|O�O�O �O�O�O�O__9_0_ B_o_f_x_�_�_�_�_ �_�_�_o5o,o>oko boto�o�o�o�o�o�o �o1(:g^p ������� � -�$�6�c�Z�l����� ��ϏƏ؏���)� � 2�_�V�h�������˟ ԟ���%��.�[� R�d�������ǯ��Я ���!��*�W�N�`� ������ÿ��̿�� ��&�S�J�\ωπ� �Ͽ϶��������� "�O�F�X߅�|ߎ߻� �����������K� B�T��x������ �������G�>�P��}�t���������  ������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<N`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz����>�y  �x�q ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^�p������q�p�x���*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p���������������$FEAT_D�EMOIN  V�� �����_INDEX����ILECOM�P [����B��8 S�ETUP2 \�BL�  �N w5_AP2�BCK 1]B	  �)����%����E �	 ���5�Y�f� �B��x/� 1/C/�g/��/�/,/ �/P/�/t/�/?�/?? �/c?u??�?(?�?�? ^?�?�?O)O�?MO�? qO O~O�O6O�OZO�O _�O%_�OI_[_�O_ _�_�_D_�_h_�_�_ 
o3o�_Wo�_{o�oo �o@o�o�ovo�o/ A�oe�o��� N�r���=�� a�s����&���͏\� 񏀏���"�K�ڏo� ������4�ɟX���� ��#���G�Y��}��@��0���ׯQ	� P�� 2� *.V1Rޯ(���*+�Q�`��W�{�e��PC��|����FR6:��"ؾg�����T   � 2����\� ��d��*.F��ϕ�	�ó����o�ߓ�STM�9���ư%�d��ψߓ�HU߻�J���f�x���GIF �A�L�-����ߑ��JPG����Lձ�n������JS�H������6���%
Ja�vaScriptt���CSe���Kֹ��v� %Casc�ading St�yle Shee�ts��j�
ARGNAME.DT'
��O�\;��[�k�|(k DISP*rUOп���� �
TPEIN�S.XML/�:�\CcCust�om Toolb�ar��	PASS�WORD���F�RS:\�� %�Passwor�d Config /c�Q/�J/�/���/ :/�/�/p/?�/)?;? �/_?�/�??$?�?H? �?l?�?O�?7O�?[O mO�?�O O�O�OVO�O zO_�O�OE_�Oi_�O b_�_._�_R_�_�_�_ o�_AoSo�_woo�o *o<o�o`o�o�o�o+ �oO�os��8 ��n��'��� ]�����z���F�ۏ j������5�ďY�k� �������B�T��x� ����C�ҟg����� ��,���P������� ��?�ί�u����(� ��Ͽ^�󿂿�)ϸ� M�ܿqσ�ϧ�6��� Z�l�ߐ�%ߴ��[� ���ߣߵ�D���h� ����3���W����� ����@����v�� ��/�A���e������ *���N���r����� =��6s�&� �\��'�K �o��4�X ���#/�G/Y/� }//�/�/B/�/f/�/ �/�/1?�/U?�/N?�? ?�?>?�?�?t?	O�? -O?O�?cO�?�OO(O��O�F�$FILE�_DGBCK 1�]���@��� < ��)
SUMMAR�Y.DG�OsLM�D:�O;_@D�iag Summ�ary<_IJ
CONSLOG1__&Q�_�_NQConsole log�_�HK	TPACCNĵ_o%o?oJUT�P Accoun�tin�_IJFR�6:IPKDMPO.ZIPsowH
�o��oKU[`Excep�tion�oyk'PMEMCHECK5o�_*_K�QMem�ory Data|L�F+l�)6qRIPE�_$6��Zs%�q Pa?cket L�_�D�L�$�	r�qST�AT���S� �%�rStat�usT��	FTP����:���Vw�Qm�ment TBD�؏� >I)E?THERNE����
q�[�NQEth�ern�p�Pfig�ura�oODDCSVRF̏��ďݟ�d��� veri?fy all���C�M.���DIF�F՟��͟b��s��d�iffd��
q��CHG01Y�@�R�篰f�z���-?��2 ݯį֯k�v������3a�H�Z�� ���ϥ�VTRNDIAG.LS��̿޿s�^q3� O�pe���q SQno�stic�weɿ)VDEV7�D�ATt�Q�c�u�g��Vis��Devisce�Ϫ�IMG7 �o����y��s�I�magߨ�UP���ES��T�FR�S:\�� �OQU�pdates L�ist �IJg�FLEXEVENQ��X�j߃�f�F� UIF Ev���B�,�s�)
PS�RBWLD.CM���sL������PP�S_ROBOWE�L��GLo�GRAPHICS4Dy��b�t��%4D� Graphic?s Fileu��A�Oɿ�rGIG����u�
YvGi�gE�ة�BN�?� )��HADO�W�����\sS�hadow Ch�ang���vb~QRCMERR��n�\s� CFG Error��tail� &����CMSGLIB��"^�o� ��T�)�ZD����/nXwZD6 ad�zHPNOTI����
/�/ZuNot�ific��H/��AGUO�/yO?�O'? P?OOt??�?�?9?�? ]?�?O�?(O�?LO^O �?�OO�O5O�O�OkO  _�O$_6_�OZ_�O~_ �__�_C_�_�_y_o �_2o�_?oho�_�oo �o�oQo�ouo
�o @�odv�)� M�����<�N� �r������7�̏[� �����&���J�ُW� �����3�ȟڟi��� ��"�4�ßX��|��� ���A�֯e����� 0���T�f�������� ��O��s��ϩ�>� Ϳb��oϘ�'ϼ�K� ���ρ�ߥ�:�L��� p��ϔߦ�5���Y��� }���$��H���l�~� ��1�����g����  �2���V���z�	��� ��?���c���
��. ��Rd����� M�q�<� `���%�I� �/�8/J/�n/ ��/!/�/�/W/�/{/ ?"?�/F?�/j?|??�?/?�?�?�$FI�LE_FRSPRT  ���0����8�MDONLY 1�]�5�0 
 ��)MD:_V�DAEXTP.Z�ZZ�?�?_OnK�6%NO Ba�ck file <9O�4S�6Pe?�O OO�O�?�O__?>_�O b_t__�_'_�_�_]_ �_�_o(o�_Lo�_po �_}o�o5o�oYo�o  �o$�oHZ�o~ ��C�g��	� 2��V��z������ ?�ԏ�u�
���.�@�~�4VISBCKH|A&C*.VDA�|����FR:\Z��ION\DATA�\v����Vision VD�B ��ŏ���'�5��Y� �j������B�ׯ� x����1���үg��� ����X���P��t��� Ϫ�?�οc�u�ϙ� (Ͻ�L�^��ς��)� ��M���q� ߂ߧ�6� ��Z�����%��I��������:LUI_�CONFIG �^�5m��� '$ h�F{�5������)�;�I���|xq�s����������� a��� $6��G l~���K�� � 2�Vhz ���G���
/ /./�R/d/v/�/�/ �/C/�/�/�/??*? �/N?`?r?�?�?�??? �?�?�?OO&O�?JO \OnO�O�O)O�O�O�O �O�O_�O4_F_X_j_ |_�_%_�_�_�_�_�_ o�_0oBoTofoxo�o !o�o�o�o�o�o�o ,>Pbt�� ������(�:� L�^�p��������ʏ ܏���$�6�H�Z� l��������Ɵ؟� ��� �2�D�V�h��� ������¯ԯ�}�
� �.�@�R�d������� ����п�y���*� <�N�`����ϖϨϺ� ����u���&�8�J� ��[߀ߒߤ߶���_� �����"�4�F���j� |������[����� ��0�B���f�x��� ������W����� ,>��bt��� �O��(:>�  xFS��$FLUI_D�ATA _�������uRESULT� 2`�� ��T�/wi�zard/gui�ded/step�s/Expert b��//+/=/O/�a/s/�/�/�*�C�ontinue �with G�ance�/�/�/?? (?:?L?^?p?�?�?�?� T-U��90 �� �?��6�9��ps�?0O BOTOfOxO�O�O�O�O �O�O�O� �_/_A_ S_e_w_�_�_�_�_�_��_�_n�?�?�?�<Frip�Oo�o �o�o�o�o�o�o! 3E_i{��� ������/�A�@S�o$on�HoAO��TimeUS/DST[������ +�=�O�a�s������'?Enabl�/˟ ݟ���%�7�I�[�Pm������T�?`{�ݯ����Æ24Ώ 3�E�W�i�{������� ÿտ翦����/�A� S�e�wωϛϭϿ��� ���ϴ�Ưد� G�~�Region�� �ߙ߽߫����������)�;�+Americasou��� �����������)�;��?�y�#߅�G�|Y��ditorL� ������#5GY�k}��+ Tou�ch Panel� �� (reco/mmen�)�� �*<N`r��U��e�w����|����accesd� ./@/R/d/v/�/�/�/�/�/�/Q|Con�nect to Network�/ (?:?L?^?p?�?�?�?��?�?�?�?Y���������!/��I�ntroduct s߆O�O�O�O�O�O�O __(_:_U^_p_�_ �_�_�_�_�_�_ oo$o6oHo e�Oeo ?O�X_�o�o�o�o '9K]o�� R_������#��5�G�Y�k�}�����h`�ooj}oߏ�o� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ쯫���Ϗ1�� X�j�|�������Ŀֿ �����0��A�f� xϊϜϮ��������� ��,�>���_�!��� E��߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~���O߱�s� ������ 2DV hz������ ��
.@Rdv ��������/ ��'/���`/r/�/�/ �/�/�/�/�/??&? 8?�\?n?�?�?�?�? �?�?�?�?O"O4O� UO/yO�OO?�O�O�O �O�O__0_B_T_f_ x_�_I?�_�_�_�_�_ oo,o>oPoboto�o EO�OiO�o�o�O (:L^p��� ����_ ��$�6� H�Z�l�~�������Ə ؏�o�o�o�/��oV� h�z�������ԟ� ��
��.��R�d�v� ��������Я���� �*��������C� ����̿޿���&� 8�J�\�nπ�?��϶� ���������"�4�F� X�j�|ߎ�M�_�q��� ������0�B�T�f� x����������� ��,�>�P�b�t��� �����������߱��� %��L^p��� ���� $�� 5Zl~���� ���/ /2/��S/ w/9�/�/�/�/�/ �/
??.?@?R?d?v? �?�/�?�?�?�?�?O O*O<ONO`OrO�OC/ �Og/�O�/�O__&_ 8_J_\_n_�_�_�_�_ �_�_�?�_o"o4oFo Xojo|o�o�o�o�o�o �O�o�O�O�oTf x������� ��,��_P�b�t��� ������Ώ����� (��oI�m��C��� ��ʟܟ� ��$�6� H�Z�l�~�=�����Ư د���� �2�D�V� h�z�9���]���ѿ�� ��
��.�@�R�d�v� �ϚϬϾ��Ϗ���� �*�<�N�`�r߄ߖ� �ߺ��ߋ�տ����#� �J�\�n����� ���������"���F� X�j�|����������� ���������� u7������ ,>Pbt3� ������// (/:/L/^/p/�/AS e�/��/ ??$?6? H?Z?l?~?�?�?�?�? ��?�?O O2ODOVO hOzO�O�O�O�O�O�/ �/�/_�/@_R_d_v_ �_�_�_�_�_�_�_o o�?)oNo`oro�o�o �o�o�o�o�o& �OG	_k-_��� �����"�4�F� X�j�|������ď֏ �����0�B�T�f� x�7��[����� ��,�>�P�b�t��� ������ί����� (�:�L�^�p������� ��ʿ��뿭��џӿ H�Z�l�~ϐϢϴ��� ������� �߯D�V� h�zߌߞ߰������� ��
��ۿ=���a�s� 7ߚ���������� �*�<�N�`�r�1ߖ� ����������& 8J\n-�w�Q� �����"4F Xj|������ ��//0/B/T/f/ x/�/�/�/�/�� �/?�>?P?b?t?�? �?�?�?�?�?�?OO �:OLO^OpO�O�O�O �O�O�O�O __�/�/ �/?i_+?�_�_�_�_ �_�_�_o o2oDoVo ho'O�o�o�o�o�o�o �o
.@Rdv 5_G_Y_�}_��� �*�<�N�`�r����� ����yoޏ����&� 8�J�\�n��������� ȟ�����4�F� X�j�|�������į֯ ����ˏ�B�T�f� x���������ҿ��� ��ٟ;���_�!��� �Ϫϼ��������� (�:�L�^�p߁ϔߦ� �������� ��$�6� H�Z�l�+ύ�Oϱ�s� ������� �2�D�V� h�z������������� ��
.@Rdv ����}���� ���<N`r�� �����//�� 8/J/\/n/�/�/�/�/ �/�/�/�/?�1?� U?g?+/�?�?�?�?�? �?�?OO0OBOTOfO %/�O�O�O�O�O�O�O __,_>_P_b_!?k? E?�_�_{?�_�_oo (o:oLo^opo�o�o�o �owO�o�o $6 HZl~���s_ �_�_���_2�D�V� h�z�������ԏ� ��
��o.�@�R�d�v� ��������П���� ����]������ ����̯ޯ���&� 8�J�\���������� ȿڿ����"�4�F� X�j�)�;�M���q��� ������0�B�T�f� xߊߜ߮�m������� ��,�>�P�b�t�� ����{ύϟ���� (�:�L�^�p������� �������� ��6 HZl~���� �����/��S �z������ �
//./@/R/d/u �/�/�/�/�/�/�/? ?*?<?N?`?�?C �?g�?�?�?OO&O 8OJO\OnO�O�O�O�O u/�O�O�O_"_4_F_ X_j_|_�_�_�_q?�_ �?�_�?�_0oBoTofo xo�o�o�o�o�o�o�o �O,>Pbt� ��������_ %��_I�[������� ��ʏ܏� ��$�6� H�Z�~�������Ɵ ؟���� �2�D�V� �_�9�����o�ԯ� ��
��.�@�R�d�v� ������k�п���� �*�<�N�`�rτϖ� ��g�����������&� 8�J�\�n߀ߒߤ߶� �������߽�"�4�F� X�j�|�������� �����������Q�� x��������������� ,>P�t� ������ (:L^�/�A�� e���� //$/6/ H/Z/l/~/�/�/a�/ �/�/�/? ?2?D?V? h?z?�?�?�?o�� �?�O.O@OROdOvO �O�O�O�O�O�O�O�/ _*_<_N_`_r_�_�_ �_�_�_�_�_o�?#o �?Go	Ono�o�o�o�o �o�o�o�o"4F Xio|����� ����0�B�T�o u�7o��[o��ҏ��� ��,�>�P�b�t��� ����iΟ����� (�:�L�^�p������� e�ǯ��믭���$�6� H�Z�l�~�������ƿ ؿ����� �2�D�V� h�zόϞϰ������� �Ϸ��ۯ=�O��v� �ߚ߬߾�������� �*�<�N��r��� �����������&� 8�J�	�S�-�w���c� ��������"4F Xj|��_��� ��0BTf x��[������ ��/,/>/P/b/t/�/ �/�/�/�/�/�/�? (?:?L?^?p?�?�?�? �?�?�?�?���� EO/lO~O�O�O�O�O �O�O�O_ _2_D_? h_z_�_�_�_�_�_�_ �_
oo.o@oRoO#O 5O�oYO�o�o�o�o *<N`r�� U_������&� 8�J�\�n�������co uo�o鏫o�"�4�F� X�j�|�������ğ֟ 蟧���0�B�T�f� x���������ү��� ���ُ;���b�t��� ������ο���� (�:�L�]�pςϔϦ� �������� ��$�6� H��i�+���O����� ������� �2�D�V� h�z���]������� ��
��.�@�R�d�v� ����Y߻�}����ߣ� *<N`r�� �������& 8J\n���� �����/��1/C/ j/|/�/�/�/�/�/ �/�/??0?B?f? x?�?�?�?�?�?�?�? OO,O>O�G/!/kO �OW/�O�O�O�O__ (_:_L_^_p_�_�_S? �_�_�_�_ oo$o6o HoZolo~o�oOO�OsO �o�o�O 2DV hz������ �_
��.�@�R�d�v� ��������Џ⏡o�o �o�o9��o`�r����� ����̟ޟ���&� 8��\�n��������� ȯگ����"�4�F� ��)���M���Ŀֿ �����0�B�T�f� xϊ�I����������� ��,�>�P�b�t߆� ��W�i�{��ߟ��� (�:�L�^�p���� ����������$�6� H�Z�l�~��������� ��������/��V hz������ �
.@Qdv �������/ /*/</��]/�/C �/�/�/�/�/??&? 8?J?\?n?�?�?Q�? �?�?�?�?O"O4OFO XOjO|O�OM/�Oq/�O �/�O__0_B_T_f_ x_�_�_�_�_�_�_�? oo,o>oPoboto�o �o�o�o�o�o�O�O %7�_^p��� ���� ��$�6� �_Z�l�~�������Ə ؏���� �2��o; _���K��ԟ� ��
��.�@�R�d�v� ��G�����Я���� �*�<�N�`�r���C� ��g���ۿ����&� 8�J�\�nπϒϤ϶� ���ϙ����"�4�F� X�j�|ߎߠ߲����� ������˿-��T�f� x������������ ��,���P�b�t��� ������������ (:����A� ���� $6 HZl~=���� ���/ /2/D/V/ h/z/�/K]o�/� �/
??.?@?R?d?v? �?�?�?�?�?��?O O*O<ONO`OrO�O�O �O�O�O�O�/�O�/#_ �/J_\_n_�_�_�_�_ �_�_�_�_o"o4oE_ Xojo|o�o�o�o�o�o �o�o0�OQ_ u7_������ ��,�>�P�b�t��� Eo����Ώ����� (�:�L�^�p���A�� eǟ��� ��$�6� H�Z�l�~�������Ư د����� �2�D�V� h�z�������¿Կ�� �����+��R�d�v� �ϚϬϾ�������� �*��N�`�r߄ߖ� �ߺ���������&� �/�	�S�}�?Ϥ�� ���������"�4�F� X�j�|�;ߠ������� ����0BTf x7��[����� ,>Pbt� �������// (/:/L/^/p/�/�/�/ �/�/����!?� H?Z?l?~?�?�?�?�? �?�?�?O O�DOVO hOzO�O�O�O�O�O�O �O
__._�/�/?s_ 5?�_�_�_�_�_�_o o*o<oNo`oro1O�o �o�o�o�o�o& 8J\n�?_Q_c_ ��_���"�4�F� X�j�|�������ď�o Տ����0�B�T�f� x���������ҟ�� ���>�P�b�t��� ������ί���� (�9�L�^�p������� ��ʿܿ� ��$�� E��i�+��Ϣϴ��� ������� �2�D�V� h�z�9��߰������� ��
��.�@�R�d�v� 5ϗ�Yϻ�}����� �*�<�N�`�r����� ����������& 8J\n���� ��������F Xj|����� ��//��B/T/f/ x/�/�/�/�/�/�/�/ ??�#�G?q?3 �?�?�?�?�?�?OO (O:OLO^OpO//�O�O �O�O�O�O __$_6_ H_Z_l_+?u?O?�_�_ �?�_�_o o2oDoVo hozo�o�o�o�o�O�o �o
.@Rdv ����}_�_�_�_ ��_<�N�`�r����� ����̏ޏ�����o 8�J�\�n��������� ȟڟ����"��� �g�)�������į֯ �����0�B�T�f� %���������ҿ��� ��,�>�P�b�t�3� E�W���{������� (�:�L�^�p߂ߔߦ� ��w����� ��$�6� H�Z�l�~������ ��������2�D�V� h�z������������� ��
-�@Rdv ������� ��9��]��� �����//&/ 8/J/\/n/-�/�/�/ �/�/�/�/?"?4?F? X?j?)�?M�?qs? �?�?OO0OBOTOfO xO�O�O�O�O/�O�O __,_>_P_b_t_�_ �_�_�_{?�_�?oo �O:oLo^opo�o�o�o �o�o�o�o �O6 HZl~���� �����_o�_;� e�'o������ԏ� ��
��.�@�R�d�# ��������П���� �*�<�N�`��i�C� ����y�ޯ���&� 8�J�\�n��������� u�ڿ����"�4�F� X�j�|ώϠϲ�q��� ����	�˯0�B�T�f� xߊߜ߮��������� �ǿ,�>�P�b�t�� ������������ ������[�߂����� �������� $6 HZ�~���� ��� 2DV h'�9�K��o��� �
//./@/R/d/v/ �/�/�/k�/�/�/? ?*?<?N?`?r?�?�? �?�?y�?��?�&O 8OJO\OnO�O�O�O�O �O�O�O�O_!O4_F_ X_j_|_�_�_�_�_�_ �_�_o�?-o�?QoO xo�o�o�o�o�o�o�o ,>Pb!_� �������� (�:�L�^�o�Ao�� eog�܏� ��$�6� H�Z�l�~�������s ؟���� �2�D�V� h�z�������o�ѯ�� ���˟.�@�R�d�v� ��������п���� ş*�<�N�`�rτϖ� �Ϻ����������� �/�Y���ߒߤ߶� ���������"�4�F� X��|�������� ������0�B�T�� ]�7߁���m������� ,>Pbt� ��i���� (:L^p��� e�w��������$/6/ H/Z/l/~/�/�/�/�/ �/�/�/� ?2?D?V? h?z?�?�?�?�?�?�? �?
O���OO/vO �O�O�O�O�O�O�O_ _*_<_N_?r_�_�_ �_�_�_�_�_oo&o 8oJo\oO-O?O�ocO �o�o�o�o"4F Xj|��__�� ����0�B�T�f� x�������moϏ�o� �o�,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ���!�� E��l�~�������ƿ ؿ���� �2�D�V� �zόϞϰ������� ��
��.�@�R��s� 5���Y�[�������� �*�<�N�`�r��� ��g���������&� 8�J�\�n�������c� ����������"4F Xj|����� ����0BTf x������� ������#/M/t/�/ �/�/�/�/�/�/?? (?:?L?p?�?�?�? �?�?�?�? OO$O6O HO/Q/+/uO�Oa/�O �O�O�O_ _2_D_V_ h_z_�_�_]?�_�_�_ �_
oo.o@oRodovo �o�oYOkO}O�O�o�O *<N`r�� ������_�&� 8�J�\�n��������� ȏڏ����o�o�oC� j�|�������ğ֟ �����0�B��f� x���������ү��� ��,�>�P��!�3�������$FMR2_GRP 1a���� �C4  B�[�	 [�߿�ܰ�E�� F@ �5W�S�ܰJ���NJk�I�'PKHu��IP�sF!��͏?�  W�S�ܰ9��<9�8�96C'6<,5����A�  �Ϲ�BH�ٳB�հ����@ӻ33�33S��۴��ܰ@UUT�'�@��8��W�>u�.�>*��<�����=[�B=����=|	<��K�<�q�=��mo���8��x	7H<8��^6�Hc7��x?�����������"��F�X���_C�FG b»T �Q����X�N�O º
F�0�� ��W�RM_�CHKTYP  ���[�ʰ̰����R{OM�_MIN�[���9����X���SSBh�c��? ݶf��[�]����^�TP__DEF_O�[��ʳ��IRCOM����$GENO�VRD_DO.��d���THR.� dzd��_ENB��{ ��RAVC��udO�Z� ����Fs  G!� �GɃ�I�C��I(i J���+���%����ʷ �QOU��j�¼������<6�i�C�;]��[�C�  D0�+��@���B����.��R SMT��k_	ΰ\����$HOSTC�h�1l¹[��\d�۰ MC[����/Z�  2�7.0� 1�/  e�/??'?9?G: �/j?|?�?�?�,Z?T3�	anonymouy �?�?	OO-O?N�/ڰRHRK�/�?�O �/�O�O�O�O_V?3_ E_W_i_�O&_�?�_�_ �_�_�_@O�_dOvOSo �_�Ojo�o�o�o�o_ �o+=`o�_�_ �����o&o8o JoL9��o]�o����� ���oɏۏ����4� j+�Y�k�}������ ��� ��T�1�C� U�g�����������ӯ ��x�>��-�?�Q�c� ����Ο���Ͽ�� ��)�;ς�_�qσ� �ϧ�ʿ ������ %�7�~�����߶ϣ� ����������Ϻ�3� E�W�i�ߍ��ϱ��� ������@�R�d�v�x� J��߉���������� ��+=`�������:$h!E�NT 1m sP!V  7 ?.c&�J �n���/�)/ �M//q/4/�/X/j/ �/�/�/�/?�/7?�/ ?m?0?�?T?�?x?�? �?�?O�?3O�?WOO {O>O�ObO�O�O�O�O �O_�OA__e_(_:_��_^_�_�_�_�ZQUICC0�_�_�_?od1@oo.o�od�2�olo~o�o!ROUTER�o�o�o�/!PCJOG�0!192�.168.0.1�0	o�SCAMPRYT�\!pu1yp��vRT�o���� !Softw�are Oper�ator Pan�el�mn��NA�ME !�
!�ROBO�v�S_�CFG 1l�	� �Au�to-start{ed'�FTP2��I�K2��V�h� z�������ԟ��� �	���@�R�d�v��� 	�������:��� )�;�M�_�&������� ��˿�p���%�7� I�[��"�4�F�ڿ�� ������!�3���W� i�{ߍߟ���D����� ����/�vψϚ�w� �ߛ��Ͽ�������� �+�=�O�a������ ����������8�J�\� n�p�]����� �����#5X �k}���� 0/D1/xU/g/ y/�/RH/�/�/�/�/ /?�/??Q?c?u?�? ���/?�?:/O )O;OMO_O&?�O�O�O �O�O�?pO__%_7_ I_[_�?�?�?t_�O�_ O�_�_o!o3o�OWo io{o�o�_�oDo�o�o��o����_ER�R n��-=vP�DUSIZ  j�`^�P�Tt>mu?WRD ?΅�Q��  guest�f�������~�SCDMNGRP 2o΅wWp��Q�`���fKL� 	�P01.05 8~�Q   �|���  ;|���  z[ ����w���*����Ť�x�������[ݏȏ���ʑPԠ������)/����D�r��ꉫ؊p"�Pl�P���Dx��dx�*���|��%�_GROU7�UpLyN��	/�\o���QUP��U�Tu� �TYà�L}?pTTP_A�UTH 1qL{� <!iPen'dan����o֢�!KAREL:q*������KC���ɯۯ��VISI?ON SET�9� ���P�>�h��f��� �������ҿ�����X�CTRL �rL}O�uſa
�aFFF9E3-���TFRS:DE�FAULT���FANUC We�b Server �ʅ�u�X���t@����1�C�U�g�;tWR�_CONFIG ;s;� ��=q�IDL_CPU_kPC���aBȠP��� BH��MIN��܅q��GNR_I�OFq{r�`Rx��NP�T_SIM_DO���STAL_oSCRN� �.��INTPMODN�TOLQ����RT�Y0����-�\�EN�BQ�-���OLN/K 1tL{�p������)�;�M���M�ASTE�%���SLAVE uL�|�RAMCACH�Ek�c�O^�O_CcFG������UOC������CMT_OPp���PzYCL�������_ASG 19v;��q
 O�r ��������&8J\W�EN�UMzsPy
��I�P����RTRY_CN��M�=�zs����Tu ������w����p/�p��P_M�EMBERS 2Yx;�l� $��X"���?�Q'W/i)��R�CA_ACC 2�y�  X�m�v 6`| �` 5�  6�i���$�&6�C�N0�/�$���b�,�$�BUF001 2�z�= l�u0  u0l�:4U�:4�:4�:4�:3�mb4b4/b4A�b4Qb4eb4vb4|�"{�"�iX:3iUj�4z�4��4��4U��4Ī4Ԫ4�4��:3j�4�4.��4Gu0�VX�j�4jk�4|�4���4��4��4��4�j�4��4�:3kbDUbD)bD9bDLbD�\bDmbD�u0�(gk�u0F��.hk�bDIDk�QDk�bD�:4�0_hg�l:4-:4U@:4P:4b:4r:4%�:4�:392$?63 :1@1ERI0ERQ0ERY0 ERa0:1h1mRq0mRy0 mR�0mR�0mR�0mR�0 mR�0�1�1:1�1�R�0 �R�0�R�0�R�0�R�0 �R�0�R�0�R�0:1�1��R@�R	@�R@t� `A�R!@�R)@�R 1@�R9@�RA@�RI@�R Q@�RY@�Ra@:1hAmb q@mby@mb�@mb�@mb��@mb�@mb�@mb�@s� �AmbI@t(�Amb�@mb�@ER�0Q�#��AER�@ ER�@ER�@ERPER	P@ERPERP:193-_ 65GSNrI2WSNrY2gS ��h3wSvry2�Svr�2 �Svr�2�S���3�S�r �2�S�r�2�S�r�2�S �r�2�S���3c�	B c��t C/c�1B?c �ABOc�QB_c�aB ocv�qBcv��B�cv� �B�cv��@v��@v��B �cv�c��C�cNr��C �cNr�B�cNrRsNr`Rs�Ԝ!��2{�Q4r�}ŋ���<��௑o�o��2�HIS�!2}� ܷ!� 2024-06�������П��� � 8�;  X
�Z=�M 9 hL!�� ���4�F�X�j� u�s�!������ί� ���(�:�L����� ��������ʿܿ� � �$�[�m�Z�l�~ϐ� �ϴ���������3�E� 2�D�V�h�zߌߞ߰� ������/��.�@� R�d�v������� �����*�<�N�`� r�������,P�������������&  Y@�� d�;+�Ic!�Ab� o�c gy������� �	-?Qc� �������/ /)/;/M/���/�/ �/�/�/�/�/??%? \/n/[?m??�?�?�? �?�?�?�?4?F?3OEO WOiO{O�O�O�O�O�O OO0O_/_A_S_e_ w_�_�_�_����5p�� ����o$o6o�� `�� `�k� !�fb)� Ao�o�o�o�O�Oo�o *<N`r� ��o�o����� &�8�J�\�n����� ��ȏڏ����"�4� F�}���|�������ğ ֟�����U�g�y� f�x���������ү� ���?�Q�>�P�b�t����������ο࿩�I_CFG 2~�[� H
Cycle Time��Busy�I�dl��minz�S�Upƾ�Read(��DowG�C� �W��Count>�	Num ������� `����P�ROG���U��P�)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,1�C�U��g�y�Tä�SDT_�ISOLC  ��Y� ���J2�3_DSP_EN�B  ��T���INC ��� c���A   ?�  �=���<#�
|���:�o ��2�D� a/�l���OB���C��O��ֆ�G�_GROUP 1큦�Qd<A*�����t�?���� `Q'�L�^��p�/�����������\�~�G_IN_A�UTO����POS�RE���KANJ?I_MASK0���DRELMON #��[�� by���������f�Ã���� d-���KCL_L NU�M��G$KEYL?OGGINGD�P�������LANGUAGE �U���DEF�AULT ��QL�G�����S�� ax�l`8T�H�  � `'0��� `; `fbK� e;���
*!(UT13:\ J/ L/Y/ k/}/�/�/�/�/�/�/��/$>(�H?�VLN�_DISP ����P�&�$�^4OCT3OL�0 aDz�����
�1GBOOK ��d4V�11�0[e%O!O3OEO�WOiKyM�TËIgF	�5)����O}����2_BUFF 2���� � `2 O�_�2��6_M�R_d_ �_�_�_�_�_�_�_�_ o3o*o<oNo`o�o�o�o�o���ADCS ������L�O���+=Oa�dIOw 2��k +�������� ����*�:�L�^� r���������ʏ܏����$�6�J�uuER/_ITM��d���� ��ǟٟ����!�3� E�W�i�{�������ï�կ�����7x�SE�VD��t�TYP����s������)�RSTe�eSCRN_FL 2��}�����/�A�0S�e�wϨ�TP{���b��=NGNAMp��E��dUPSf0SGI��2�����_LOAD��G �%��%PLACE_TORN �1߬6MAXUALcRMb2�@���9
K���_PR��2 � �3�AK�Ci0���qO=_'X�Ӭ�P �2��; �*V	Z����
* ��� 4��*��'�`�	xN� ��z��������� ��1�C�&�g�R���n� ����������	�� ?*cFX��� ����; 0q\����� ��/�/I/4/m/ X/�/�/�/�/�/�/�/ �/!??E?0?i?{?^? �?�?�?�?�?�?�?O OAOSO6OwObO�OD��DBGDEF ���գѢѤO�@_L?DXDISA�����ssMEMO_AP���E ?��
 �A�H$_6_H_Z_�l_~_�_�_K�FRQ_CFG ���m�CA �G@��S�@<��d%�\o�_t�P�Ґ���ԯ*Z`/\b **:eb�DXojho �F�o�o�o�o�o�o ;�O��dZ�U�y|��z,(9�Mt ���1��B�g�N� ��r��������̏	����?�A�ISC 31���K` ��O�� ���O���O֟����K��]�_MSTR ��3��SCD 1�]��l��{� ����دïկ���2� �V�A�z�e������� Կ�������@�+� =�v�aϚυϾϩ��� ������<�'�`�K� ��oߨߓߥ������ ��&��J�5�Z��k� ������������� �F�1�j�U���y��� ����������0�T?x�MK�Q�,��Q�$MLT�ARM�R�?g� ~s�@��>�@METPU�@l���4�NDSP?_ADCOL�@�!CMNT7 �*FNSW(FS�TLIxi%� �,����Q��*_POSCF�b�PRPMV�STv51�,� 4�R#�
g!|qg%w/�' c/�/�/�/�/�/�/? �/?G?)?;?}?_?q?��?�?�?�?�1*SI�NG_CHK  }{$MODA�S��e���#EDE�V 	�J	M�C:WLHSIZE��Ml �#ETASK� %�J%$12�3456789 ��O�E!GTRIG ;1�,� l�Eo�#_�y_S_�}�FYP�A�u9D"CEM_�INF 1�?k�`)AT&F�V0E0X_�])��QE0V1&A3�&B1&D2&S0&C1S0=�])ATZ�_#o
d�H'oOo�QC_wohA�o�obo�o�o�o  �_&�_�_�_o�3o ��o���o��"� 4��X���AS e֏���C�0�� �f�!���q�����s� 䟗�����͏>��b� ��s���K���w��� ٯ�ɟ۟L����#� ����Y�ʿ���� $�߿H�/�l�~�1��� U�g�y����ϯ� �2� i�V�	�z�5ߋ߰ߗ�|��PONITOR��G ?kK   	EXEC1o��2�3�4�5���@�7�8�9o����(� ��4��@��L��X �d��p��|��2���2��2��2��2���2��2��2��2���2��3��3��3�(�#AR_GRP_�SV 1��[ �(�1?��>����	>��>-��׿�8��3�RM�A_DsҔN~��ION_DB-@��1Ml  �J� w� xJD"�� -�/��FH���N   22V�/ .yJE-u�d1}E���)P�L_NAME �!�E� �!D�efault P�ersonali�ty (from� FD)b (RR�2�� 1�L��XL�p�X  d�-?Qc u������� //)/;/M/_/q/�/�/�/EC2)�/�/�/ ??,?>?P?b?t?EB<�/�?�?�?�?�?�?�
OO.O@OROdO��6�?�N
�O�O�P�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_�O�O2oDoVoho zo�o�o�o�o�o�o�o 
.@o!ov� ���������*�<�N�`�r������ Fs  GT?�G�M����  �ÏՍ�d �������(�6��� ���
 �m�~�h����� ������ğ֟ �����:���
�]�m����	`������|į��:�oA������ A�  /���P���� r�������^�˿ݿȿ���%��R�� 1��	X ��, �� ��� a� �@D�  t�?��z�`�?� |��A/���t�S��;�	�l��	 ��xJ���x��� �� �<�@����� ��·�K��K ��K�=*�J���J���J9���
�ԏC߷�@�t��@{S�\��(�Ehє��.��Iߑ��ڌ����T;f�ґ�$��3��´  �@���>�Թ�$�  >�����ӧf  � ��x`���� R� ���Ǌ���� �  { � @T�����  �  �l�ϊ��-�	'� � ���I� � � �<�+�:������È=��ͨ��0Ӂ��N �[��n @���f����f�k���,�av�  '��Yэ��@2��@�0�@�Ш���C��C>b C��\C����:��G�@B���
� ����� )�Bb $/�!��L�Dz�o�ߓ�~��0��( �� -���������!9��D�  9�恀?��ffG�*<� !}�q�1�89�B�>��bp��(�(9��P��	������>�?��9�x9��W�<
6b<���;܍�<����<���<�^���I/��A�{���fÌ�,�?fff�?_�?&� T�@��.�"�J<?�;\��"N\�6��� �!��(�|��/z��/j' ��[0??T???x?c? �?�?�?�?�?�?6��%F���?2O�?VO�/�wO�)IO�OEHG@� G@09�G�� G}ଙO�O�O_�	_B_-_f_Q_BL
9�B��Aw_[_�_b� �_�[�_��mO3o�OZo��_~o�o�o�o���bs��PV( @|po 	lo-*cU�ߡ!A���r59�CP�xLo�}?�����#��6��W9����6�Cv�q�CH3� j�t����q������|^(hA� ��ALffA]���?�$�?���;�°u�æ��)�	ff��?C�#�
����g\)�"�33C��
�����<��؎G�B����L�B��s�����	";�H�ۚG���!G��WI�YE���C��+�8�I۪�I�5�HgM�G�3E��R�C�j=x�
�p�I���G��f�IV=�E<YD�C<�ݟȟ�� ��7�"�[�F��j��� ����ٯį���!�� E�0�i�T�f�����ÿ ���ҿ����A�,� e�Pω�tϭϘ��ϼ� �����+��O�:�s� ^߃ߩߔ��߸����� � �9�$�6�o�Z�� ~������������ 5� �Y�D�}�h����� ����������
C:.(䁳��/"����<��xt��q3�8��<��q4Mgu����q�VwQ�
4p�+4�]$ $dR�v���u%PD"P��Q�_/�Z/=/(/a/L+R�g/n/�/�/�/�/�/  %��/�/+??O? :?s?/�_�?�?�?�;�?�?O�? OFO4O�rLO^O�O�O�O��O�O�J  2 {Fs�wGT�V�M�uBO�|r�pp�C��S@�R_�p�oy_�_^_�_o 6\!�WɃ�_o�o(o�z?���@U@�z�D�p�p�k1�p�~
  6o�o�o�o�o�o�o );M_q�ڊ�sa ����D���$MR_CA�BLE 2��O ]��T�	LaMa?�PMaLb�pK�Z��&P�C�p�?aO4>�B����?a��}?`?aE)~�?f��v��l  ��&Pļv�wdN�{0���$P ��cF �%� 6�H�XT���6P?`C$�ČZ��n��k&�g�������� �ɾ&P��C���=�u��ǌ�j�?`z�Z<v։��s 9��T�,�>���b��� ����Ɵ��Ο3�.�� P�(�:���^�����#?`������<h�pH�Z�l�<h*���** �sOM }��y���B?b�6=%% 23�45678901�ɿ۵ ƿ���?`�h?`AQ!�?a
��z�not segnt ���W��TESTFE�CSALG� egD;jAQd��ga%�
���@��?d�r���������� 9U�D1:\main�tenancesG.xmS�.�@�vj��DEFAU�LT�\�rGRP {2���  pld��G?e  �%1�st mecha�nical ch'eck�?aՀ��#������E��Z��(�:�L�^�?b��c�ontrolleAr�Ԍ��߰��D������ ��$�s�M��L�?b"8b���v��B�����������/�C}�a�6����dv���s��C��ge��. b?attery�&��E	S(:L^�p�	|�duiz�awblet  D��"��R����/"/4/s��g�reas�>gf�Br#-?`|!�/�E�@�/�/�/�/�/s�
��oi,�g/y/�/��/t?�?�?�?�?s�H�
�?f�W��1<?`AO�E
c?8OJO\OnO�O�t��?O��'O�O_ _2_D_s��OverhaulE��L��R x?`�Q�_���O�_�_�_�_o?`$�_0o����_o �_�o�o�o�o�o o�o?oQocoJ\ n���o�) ��"�4�F���|� �k��ď֏���� [�0�B���f������� ����ҟ!���E�W�,� {�P�b�t�����矼� ���A��(�:�L� ^�����ѯ㯸��ܿ � ��$�s�Hϗ��� ~�Ϳ�ϴ�������9� �]�o�Dߓ�h�zߌ� �߰�����#�5�G��� .�@�R�d�v��ߚ��� ���������*�y� ��`���O�������� ����?�&u�J�� n�����) ;_4FXj| ����%�/ /0/B/�f/���/ ��/�/�/�/?W/,? {/�/b?�/�?�?�?�? �??�?A?S?(Ow?LO ^OpO�O�O�?�OOO +O�O_$_6_H_Z_�O ~_�O�O�O�_�_�_�_po o�PeR	 T"o Ooaoso�_�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
���  ��Q?�w  @eQ �o W�i�{�eVC�����̟�bX*�**  �Q�V��� �2�D��ph�z��������_ �S������կ7� I�[�����ɯ/���ǿ ٿ#���!�3�}��� ��{ύϟ��s����� ��C�U�g��S�e�w߀9ߛ߭߿�	��eU�eQ�$MR_HI_ST 2��U��� 
 \jR$ �23456789C01*�2����)�9c_���R��a_�� �������=�O�a�� *�x�����r����� ��9��]o&� J�����# �G�k}4�Z��SKCFMAPw  �U�)���Z���ONREL  �����лEX_CFENB'
���!FNC$/$JOGOVLIM'qd�m �KEY'�p%y%_PANp(�"�"�RUN`,�p%�SFSP�DTYPD(%�S�IGN/$T1M�OTb/!�_C�E_GRP 1��U�"�:`��n? Z[?�?�؆?�?~?�? �?�?!O�?EO�?:O{O 2O�O�OhO�O�O�O_ �O/_�O(_e__�_�_ �_�_v_�_�_�_o����QZ_EDIT�4��#TCOM_�CFG 1���'%to�o�o 
Ua_/ARC_!"��O)�T_MN_MOD�E6�Lj_SP�L�o2&UAP_C�PL�o3$NOCH�ECK ?� � Rdv ����������*�<�N�`��NO_WAIT_L 7lJg50NT]a����UZ��_ERR&?12���ф��	� �-����R�d����`�O����| 6`��
aB���ƒA�&����<���I�@�,W<� �� ?��j�ϟj����قP�ARAMႳ��N�oR�=��o��� = e���� ��گ�ȯ��"�4��0X�j�F�<�蜿���A�ҿ�"ODRDS�P�c6/(OFFS?ET_CAR@`�o��DIS��S_�A�`ARK7KiO�PEN_FILE�4�1�aKf�`OPT?ION_IO�/�!���M_PRG %�%$*����h��WOT��E7�O����Z��  %��"�÷"�G	 �W"�Z����RG_DS�BL  ���ˊ���RIENTkTO ZC����A �U�`IM�_D���O��V~�LCT ����Gbԛa�Zd��_�PEX�`7�*�RA-T�g d/%*���UP ���{��������������/$PAL�������_POS_CHU��7����2>3�L��XL�p��$�ÿU�g�y��� ������������	 -?Qcu����Y2C���" 4FXj|�� ���� //$/6/@H/Z/l/~/�Y�� �.��/�/ςP�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO�/ �/LO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_)O;O�_�_�_�_�_ �_�_o o2oDoVoho�zo�o�o�_<�� �o�m ���(�"{ BPw�m�m���~�jw8��w���� ��2�T��p��w���H��t	`���̏ޏ��:�o������ �2��pA�   I��j�`������ ���џ���@���#�)�Or�1����� 8�>��, �\Ԡ�~� @D�  ��?���~�?� ���!�D������%G� � ;�	l��	 ��x�J젌����� ��<� ��� ���2�H(��H�3k7HSM5G��22G���GN�3%�R��oR�d��2�Cf��a��{���������/��3��-¸��4��>����𚿬���3�A�q�½{q�!ª��ֱ� "�(«�p=�2����� ��_{  @�Њ��_�  ��Њ��2���.�	'� �� ��I� ��  �V�,�=�������˖ß���  �y��n @"��]�<߭�"������-�N�Д߇  '�Ь�w�ӰC>��C��\C߰���Ϲ��ߤ!���@%�4���/��2�~�B��B�I�;�)�j客z+���쿱����������( �� -��#�������!�]�9�|�  q�?�ffaH�Z��� ������"��8� ����>�|P$��}�(� ��P��������\�?���� x� ���<
6�b<߈;܍��<�ê<���<�^�*�gv�A)ۙ�脣��F��?fff?}�?&�� ��@�.���J<?�\��N\��)������� ����ޤy�N9 r]������ �/&/�J/5/n/��	g/�/c(G@� G@0i�G�� G}���/??<?�'?`?K?�?o?BL
i�B��A�?y?�?|� �?K�?ů�/QO�/xO��?�O�O�O�Om��bs��n�t @|�O '_�OK_6_H_�_lS��!A��RS�i�Cn_�_xj_0O�]?��o�oAo,où�Wi����ToC���`CH�Qo>Jd�`a�a@�Iܚ>(hA�� �ALffA�]��?�$�?����ź°u��æ�)�	ff���C�#�
ܢopg\)��3�3C�
������<��nG��B���L��B�s�����	0źH����G��!G���WIYE����C�+�½I�۪I�5�H�gMG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo�� �
��U�@�y�d��� ������я����� ?�*�c�N���r����� ���̟��)��9� _�J���n�����˯�� �گ�%��I�4�m� X���|���ǿ���ֿ ���3��W�B�Tύ� xϱϜ���������	� /��S�>�w�bߛ߆� �ߪ߼�������=��(�a�L�(q���)����Z�������a3�8�������a4Mgux�����a�VwQ��(�4p�+4�]B�B���p�����������UPbP���Q O%x�1[FjR�������  C���I 4mX�8
O������.//>/d/R/�Rj/|/�/�/�/�/�/:  2� Fs�gGT]�&6�M�eBmpX�R�P�aC��3@�_ p?�?�?�?�?�?�=�S�OO)O;OMO�c�?���@@�jJ��`�`�1�`�^
 TO�O�O �O�O�O_#_5_G_Y_�k_}_�_�_�j�A �����D��$�PARAM_ME�NU ?B���  �DEFPULS�E�[	WAIT�TMOUTkR�CVo SH�ELL_WRK.�$CUR_STY�L`DlOPT�Z1ZoPTBooibC�?oR_DECSN `���l�o�o�o &OJ\n������QSSREL_ID  >��
1��uUSE_P�ROG %�Z%8�@��sCCR` ��
1�SS�_HOST7 !�Z!X����M�T _���x�������L�_TIME�b �h��PGDE�BUG�p�[�sGI�NP_FLMSK��E�T� V�G�PG�Ar� 5��?��CyHS�D�TYPE�\�0��
�3�.� @�R�{�v�����ï�� Я����*�S�N� `�r����������޿ ��+�&�8�J�s�n���ϒϻ�G�WORD� ?	�[
 	�PR2��MA9I�`�SU�a��cTEԀ���	Sd�COL��C߸��L� C�~��h�d*�TRACE�CTL 1�B���Q ��b c'��0�ށ�_DT Q�B������D � ��|A��	��
���������Հ1�@�@����P�A�@������T ���������U��OF�ON�OV�UO^�Of�On�Ov�Qx�S0z�x�x�� z�x�x�@��U�^��f��n��F�U�N������&�����6��>��Ң��&���7��>�Ӫ����&�����*6��>�������:W�� ��	!Q������&����U�6��>�Ѯ�Ѷ��-?Qc	������J��������V���o��'���O��O�6�O>�O��O��O���O��O��O�O �M�_�����%�7� I�[�m������� ��������3�E�O i�{�������k��T�#'3�.4�64�nQЎ%�O�O� �+=�*���� (O:OLO^OpO�O�O�O �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� P�$Or���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~�f������  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o�o�o�o�a�$PG�TRACELEN�  �a  �_��`��f�_UP �����q'pq� p�a_CFG M�u	s�a p�LtLtfqwpqz�  �qu4rD�EFSPD ��?|�ap��`H�_CONFIG s�us �`��`d�t��b ��a�qP�t�q��`���`IN7pTRL' �?}_q8�u��PE�u��w��qLt�qqv�`LI�D8s�?}	v�LL�B 1��y k��B�pB4Ńqv �އ؏	��s << �a?��'���A� o�U�w�������۟���ӟ��#�	�+�Y�v� 񂍯����ï
���������/�u�GRP �1ƪ��a@俼j��hs�aA��
D�� D�@� Cŀ @�٭^�t�q�����q�p���.� ���FȾ´���ʻB� )�	���?�)�c��a�>��>�,���Ϻ��ζ� =49X=H�9��
��� �@�+�d�O���s߬��o߼�����  Dz���`
��8���H� n�Y��}������� ������4��X�C�|����)��
V7.10beta1Xv A�������!�����?!G��>\=y��#��{33A!�ߚ@��͵��8�wA��@� A�s�@Ls���� ��"4FXLsA�pLry�ā���_��@l��@ë33q�`s��k���Anff�a���ھ��)�x�� �ar�T� n�t����	t��KNOW_M  �|uGvz�SV ��z�r�&�� ��>/�/G/�aԤ�y�MM���{ ����	^u (�l+/�/',_t@oXLs�����@���%�"4�.�N�z�MRM��|-T�U�y�c?u;eOADBANFWD~�x�STM�1 1��y�4Ga�rra_B�2Se�m��?~s�;CEo�2��O�7�3�Antena_F?ull @��VO De�qH��^OpO�O�O �O�O�O�O!_ __W_ 6_H_�_l_~_�_�b�7�2�<�!4�_  �#<�_�_N�3�_�_
oo�749oKo]ooo��75�o�o�o�o�76 �o�o�772DVh�78����V�7MA�0��s�wwOVLD  ��{�/a�2PAR?NUM  �;]���u�SCH*� �8�
����ω�3�U�PD��[�ܵ+�wu_CMP_r -��0��'�5C�ER_C;HKQ����1�"e�N�`�RS>0�?G�'_MO�?_��#u�_RES_G�0��{
Ϳ@�3�d�W� ��{��������կ����*�����P� �O��8`l������ �`��ʿϿ��`�	� ��1p)�H�M���p hχό���p�������V 1��5�1�!�@`y�ŒTHR_INR>0/�Z"z�5d:�MASSGߛ Z[�MNF�y�M�ON_QUEUE� ��5�6Ӑ~  U#tNH�U��N������END������EXE�����BE�������OPTIO�������PROGR�AM %��%���߰���TASK�_I,�>�OCFG� ά�]�����D�ATAu#������	�"2 �O=���`�r�����:�� ������������� ~
1C�U�INFOu#� ���Ԕ$���� ��
.@Rd v��������/as x� � �;���ȀK_���8��S&ENB-�b-�&q�&2�/�(G��2��b+ X,	�	��=����/�'�@��P4$�0���99)�N'_EDIT ���W?i?��WERFL�-ӱ3�RGADJ �F:AN�5?Ӑ�5W��6��]!֐���?�  BzD�WӐ<1Ӑ�%�`%O�8;��50!2��7֊	H��l0��,�BP�0�@\�0�M*�@/�B **:�B�O�F�O2��D��A�ЎO�@@O	_,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_ �_o�_o�_�_
o�o .o�ojodovo�o�o�o �o�o�o\XB< N�r����4� �0���&���J��� ������������ ��x�"�t�^�X�j�� ����ʟğ֟P���L� 6�0�B���f������� ��(�ү$������ >���z�t��� Ϫ��� ���l��h�R�L�^�DX	����1���"���t$ :�L���o�
ߓߥ��7PREOF ��:�0�0�
�5IORITY�X�M6��1MPDSaPV�:
B �UT��|�C�6ODUCT���F:��NFOG[@_TG�0��J:?��HIBIT_DO��8��TOENT �1�F; (!?AF_INE*���~��!tcp��>�!ud��8�?!icm'��N�?�XY�3�F<��1)� �A�����0����������� ' ]D�h�@�����*>��3��9
BOTf�3�>�80�F�G/��LC��4�;LFJA~B,  ��ЀF!//%/7/�5�F�Z�w/�/�/�/�3�&ENHANCOE �2FBAH+Ad�?�%;��������Ӓ1�1PORT�_NUM+��0����1_CART�RE�@��q�SK�STA*��SLGmS������C��Unothing?�?OO�۶0TEMP �N��"O�E�0_a_seiban|߅Ox� �O�O�O�O�O_�O'_ _K_6_H_�_l_�_�_ �_�_�_�_�_#ooGo 2okoVo�ozo�o�o�o �o�o�o1U@ e�v����� ����Q�<�u�.I�VERSI	�L���� disa�ble'2*KSAV�E �N�	2670H771|�	h��!�/��9��:� 	^�4�ϐ����e��͟ߟ������9�D�C-Å_�y� 1�������ő����Ǻ�URGE� B��r�WFϠ��-��9�W�����l:WRUP�_DELAY ��=n�WR_HOT %��7��/p���R_NORMA�LO�V�_�����SE�MI��������QS�KIPo��97��x f�=�b�a�sυ�H��� ���ø��������&� �J�\�n�4�Fߤߒ� �����߲���� �F� X�j�0��|������ ������0�B�T���x�f���������ãR�BTIF�5���C_VTMOU�7�5����DCRo��� М�A�y�"C��C���>�.}>Ą;݆H����/t�ž���˾,̹k��HϘ�� <
�6b<߈;����>u.�>*?��<��ǪP0���2DV hz��������,GRDIO_T?YPE  v���/ED� T_CF�G ��-�BHf]�EP)�2��+7 ���B�u �/ �*��/�?�/%?= �/V?�}?�Ϟ?���? �?�?�?�?O
O@O*G l?qO��8O�O�O�O�O �O�O�O�O_<_^Oc_ �O�__�_�_�_�_�_ o�_&oH_Mol_o�o o�o�o�o�o�o�o�o "DoIho*j� ������.3� E��f� ���x����� ���ҏ�*�/�N�� b�P���t�����Ο���ޟ�:�+���R'INOT 2�R��!��G;� i�{��"�<��8f�0 ��ӫ ������M�;� q�W�������˿��� տ�%��I�7�m�� eϣϑ��ϵ������� !��E�3�i�{�aߟ� ���߱����������A���EFPOS1� 1�!)  x���n#����� ��������/��S� ��w����6�����l� ������=O���� 6���V�z � 9�]�� ��Rd���#/ �G/�k//h/�/</ �/`/�/�/??�/�/ ?g?R?�?&?�?J?�? n?�?	O�?-O�?QO�? uO�O"O4OnO�O�O�O �O_�O;_�O8_q__ �_0_�_T_�_�_�_�_ �_7o"o[o�_oo�o >o�o�oto�o�o!�o EW�o>��� ^�����A�� e� ���$�����Z�l� ����+�ƏO��s� �p���D�͟h�񟌟 �'�ԟ�o�Z��� .���R�ۯv�د��� 5�ЯY���}���*�<� v�׿¿����Ϻ�C��޿@�y��e�2 1�q��-�g�����	� �-���Q���N߇�"� ��F���j��ߎߠ߲� ��M�8�q���0�� T��������7��� [�����T������� t�����!��W�� {�:�^p� �A�e � $��Z�~/� +/���$/�/p/�/ D/�/h/�/�/�/'?�/ K?�/o?
?�?.?@?R? �?�?�?O�?5O�?YO �?VO�O*O�ONO�OrO �O�O�O�O�OU_@_y_ _�_8_�_\_�_�_�_ o�_?o�_co�_o"o \o�o�o�o|o�o) �o&_�o��B �fx��%��I� �m����,���Ǐb� 돆����3�Ώ��� ,���x���L�՟p��� ����/�ʟS��w��x���ϓ�3 1�� H�Z������6�<�Z� ��~��{���O�ؿs� ���� ϻ�Ϳ߿�z� eϞ�9���]��ρ��� ߷�@���d��ψ�#� 5�G߁�������*� ��N���K����C� ��g��������J� 5�n�	���-���Q��� ������4��X�� Q���q� ��T�x �7�[m�/ />/�b/��/!/�/ �/W/�/{/?�/(?�/ �/�/!?�?m?�?A?�? e?�?�?�?$O�?HO�? lOO�O+O=OOO�O�O �O_�O2_�OV_�OS_ �_'_�_K_�_o_�_�_ �_�_�_Ro=ovoo�o 5o�oYo�o�o�o�o <�o`�oY� ��y��&��#� \�������?�ȏ����4 1�˯u��� ��?�*�c�i���"��� F����|����)�ğ M�����F�����˯ f�﯊�����I�� m����,���P�b�t� �����3�οW��{� �xϱ�L���p��ϔ� ߸������w�bߛ� 6߿�Z���~����� =���a��߅� �2�D� ~��������'���K� ��H������@���d� ����������G2k �*�N��� �1�U� N���n��/ �/Q/�u//�/4/ �/X/j/|/�/??;? �/_?�/�??�?�?T? �?x?O�?%O�?�?�? OOjO�O>O�ObO�O �O�O!_�OE_�Oi__ �_(_:_L_�_�_�_o �_/o�_So�_Po�o$o��oHo�olo�oۏ�5 1����o�o�ol W��o�O�s� ��2��V��z�� '�9�s�ԏ������� ��@�ۏ=�v����5� ��Y��}�����۟<� '�`��������C��� ޯy����&���J�� ��	�C�����ȿc�� ��ϫ��F��j�� ��)ϲ�M�_�qϫ�� ��0���T���x��u� ��I���m��ߑ��� �����t�_��3�� W���{������:��� ^�����/�A�{��� �� ��$��H��E ~�=�a�� ���D/h� '�K���
/� ./�R/��/K/�/ �/�/k/�/�/?�/? N?�/r??�?1?�?U? g?y?�?O�?8O�?\O �?�OO}O�OQO�OuO��O�O"_t6 1�%�O�O_�_�_�_ �O�_|_o�_o;o�_ _o�_�oo�oBoTofo �o�o%�oI�om j�>�b�� �����i�T��� (���L�Տp�ҏ��� /�ʏS��w��$�6� p�џ���������=� ؟:�s����2���V� ߯z�����د9�$�]� �������@���ۿv� ����#Ͼ�G����� @ϡό���`��τ�� ��
�C���g�ߋ�&� ��J�\�nߨ�	���-� ��Q���u��r��F� ��j����������� �q�\���0���T��� x�����7��[�� ,>x��� �!�E�B{ �:�^���� �A/,/e/ /�/$/�/ H/�/�/~/?�/+?�/xO?5_GT7 1�R_ �/?H?�?�?�?�/O �?2O�?/OhOO�O'O �OKO�OoO�O�O�O._ _R_�Ov__�_5_�_ �_k_�_�_o�_<o�_ �_�_5o�o�o�oUo�o yo�o�o8�o\�o ��?Qc�� �"��F��j��g� ��;�ď_�菃���� ��ˏ�f�Q���%��� I�ҟm�ϟ���,�ǟ P��t��!�3�m�ί ��򯍯���:�կ7� p����/���S�ܿw� ����տ6�!�Z���~� Ϣ�=ϟ���s��ϗ�  ߻�D������=ߞ� ����]��߁�
��� @���d��߈�#��G� Y�k�����*���N� ��r��o���C���g� ����������n Y�-�Q�u� �4�X�|b?t48 1�?); u��/;/�_/ �\/�/0/�/T/�/x/ ?�/�/�/�/[?F?? ?�?>?�?b?�?�?�? !O�?EO�?iOOO(O bO�O�O�O�O_�O/_ �O,_e_ _�_$_�_H_ �_l_~_�_�_+ooOo �_soo�o2o�o�oho �o�o�o9�o�o�o 2�~�R�v� ��5��Y��}�� ��<�N�`������� ��C�ޏg��d���8� ��\�埀�	�����ȟ �c�N���"���F�ϯ j�̯���)�įM�� q���0�j�˿��� ��Ϯ�7�ҿ4�m�� ��,ϵ�P���tφϘ� ��3��W���{�ߟ� :ߜ���p��ߔ��� A����� �:���� Z���~�����=���a���� �����M�ASK 1���������XNO�  ���� MO�TE    �N_CFG ��Y����PL_RGANGUP���OWER ���� �A��*S�YSTEM*P�V9.3044 ��1/9/2020� A �g ����RESTART�_T   , �$FLAG� �$DSB_SIG�NAL� $U�P_CND4P���RS232r� � $COM�MENT �$DEVICEU�SE4PEEC$�PARITY4O�PBITS4FL�OWCONTRO~3TIMEOUe�6CU�M4AU�XT��5INTE�RFACsTAT}U���K�CH t �$OLD_yC�_SW 'FR�EEFROMSI�Z �ARGET�_DIR 	�$UPDT_MA�P"� TSK_E;NB"EXP:*#�!jFAUL E�V!�RV_DA�TA�  �$n E�   	�$VALU�! �	j&GRP_ �  {!A � 2 �SC�R	� �$�ITP_�" �$NUM� OUP�� �#TOT_AXܕ�#DSP�&JO�GLI�FINE�_PCd�OND��%$UM�K�5 _MIR1!4PvP TN?8APL"G0_EXb0<$�!� �814�!PGw6BR�KH�;&NC� I�S �  �2TYQP� �2�"P+ Ds<�#;0BSOC�&R �N�5DUMMY1�64�"SV_CO�DE_OP�SF�SPD_OVRD��2^LDB3OmRGTP; LEF�F�0<G� OV5S�FTJRUNWC!S�FpF5%3UFRA��JTO�LCHD�LY7RECOVD'� WS* �0�EF0RO��10_p@�   @��S� NVERT"O�FS�@C� "FW�D8A�D4A�1ENAYBZ6�0TR3$1�_`1FDO[6MB�_CM�!FPB� B�L_M��!2hRnQ2xCV�"' } �#PBGiW|8AMz3\P���U�B�__M�P�Mx� �1�AT$CA� ��PD�2�PHBK�+!:&aIO�4 �eIDX+bPPA j?a$iOd7e�U7a�CDVC_DBG"��a;!&�`�B5�e1Ƞj�S�e3�f�@AT�IO� ���AU0�c� �S�AB
0Y.#0�D��X!� �_�:&SUBCPyU%0SIN_RS�T, 1N|�S�T!��1$HW_C1��"]q.`�v�Q$A�T! � �$UNI�T�4�p�pATT�RI= �r0CYC=L3NECA�bL3�FLTR_2_F�I9a7�c,!LP�;CHK_�SCmT>3F_�wF_�|�8��zFS+�R�rCHAGp�y��R�x�RSD�@'�1E#&v7`_T�XPRO�`�@S�EMPER_D0�3Tf�]p� f���P�DIAG;%R�AILAC�c4rMF� LO�0�A�65�"PS�"�2 -`�e�SkPR�`S.  ��W�Ctaf	�CFU�NC�2�RINS_T.!(�w��&� S_� �0�P��8 	d��WARL0b?CBLCUR��єaAʛ�q͘ƘDA�00���ѓʕLD @�,a3��!��8�3�T�ID�S��!� $C�E_RIA !5AFDpPC~��@���T2 �C9#�b{QO�I�pCVDF_LE���#0(!�LM�SF}A�@HRDYOL1	PRG8�H��>1(|�ҥMULSE t=#Sw3��$JJ�J6BKGFKFAN_�ALMLV3R�W{RNY�HARD�0$+&_P "��2Q��d�!�5_�@:&AU��Rk��TO_SBRvb��� ƺ�pvc��޳MPINF�@p�q�)���REG'd�~0V) 0R�C�1DA3L_ \2FL�u�2$MԐ(�#S��P�� `�g�CMt`NF�qsONIP�q5p�IPP �9a$Y��! ��"�!� ��o3EGP��#@��AR� �c�52������|5AXE�'ROBn�*RED�&WR�@2�1_=��3SY�0�t�0_�Si�WRI�@�ƅpST�#��0*@� �q	���3��� �B� �A��3�D�PO�TO�� �@AR�Y�#��!��d�!1F�I�0�$LIN]K��GTH�B ST_���A��6�"N/�XYZ+"9�7G�'OFF�@�.�"�%��B� l����A3$ ��FI�p���h4�4l��$_Jd��"(B�,a������8@�"q������C�k6DUR��94�TURT�XZ�N����1Xx��P��FL/�@`s��l�P��30�"^Q 1� K
0	M:$�53]q7�SuD�Sw#ORQɆ�!��P���Q7��0O[�ND��=#�!#�1OVE8��M���R�� R��Q!P.!P! OAN}q	�R���� 990� �brJ9V`����v�!ER1
��	8�E�@n D�	A��p�嘕Ă���v�AX�C�"� �`�q�s�� �0~3�~F�~e�~�~E�~1��~Ҡ {Ҡ�Ҡ�Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�Ҡx�!)DEBU}s$x���삼!R*�CAB�a8A2V`|r 
�"�c���% �Q7�7�173�7 F�7e�7�7E�p������LAB��q��yp�cGRO�p4��}��PB_ҁ  ��̓��ð�6�1���5���6AND��8p �a3���-G �Q�����AH�PH�p2�NT8d��Cs@VEL؁��}A��F�SERV9Es@�� $����mA!�!�@POR }�KP�иA���@���	  $�BTRQ�
�CH��@
�G��2	�Eb��?_  lb��QN�ERR��RI�P8�@�FQTOQ�� AL�}��YVĀG�Ea%�\���BRE�  ,�A�EP�
�RA�Q 2' d�R7c�U�@7 ��$F ׂl��m d�COC���P  8[C�OUNT���@��F�ZN_CFG�A# 4�p%��rT\zs �a�#`pJp b��(a��/ �� MGp+�����`�OGp�eFAq����cX8еk�i�oQ��'ѴDp8�P~z��SHELA�~-b 5���B_BAS\RS)R$�`�2�S��L�R!p1�W!p2Dz3DzU4Dz5Dz6Dz7Dz98�WqROO���P��1�NL�� �AB��C
�"pACK�&I%N�PT+�W�U��	�k��y_PU8�~�|�OU�CP��%�s�V�l���YTPFWD�_KARKQ-�:PR�E�D�P����QUE$�Ā9 )���~���IU��#s/���@�/�SEM1ǆ1��A�aSTY�tSO����DI�q��Qc���X��_TM9�M�ANRQ �/�EN�D��$KEYSWITCH2�G�����HE)�BEATmMz�PE��LEJR(���0x�UF�F��G��S�DO_HOM���Oz��pEFPAR��SbJі��uC���O��7P�QOV_Mx��}�c�IOCM�d��1�� uHK��G D,�&�a`U2R�M��a�r +�FO;RC*�WAR���OM��  @��$�㰰U��P�1(��g���3��4�1�B*�POW�Lz��R%�OUNLO�0T��ED��  �S�NP��S.b 0�N�ADDa`z�$�SIZ*�$VA��0�UMULTIP��r���Az� � $��ƒ$���SQc�1CFPv�OFRIFr�PSw�؉�ʔf�NF#�ODBUx�R@w������F��:�IAh����������S"p�� �3  �cRTE��.�SGL.�T�x��&C`Gõ3a�/�ST�MT��`�P����ByW9 0�SHOWh�nqBANt�TPo����E������@V�_Gsb �$�PC�0�PoFBZv�P��SP��A�p�����D��rbw� �+QA002D .ҝ�6ק�6ױ�6׻��6�54�64�74�8*4�94�A4�B4و� 6ׇ17�}�6�F4�  ��@�����Z����t�U1��1��1��1��U1��1��1��1��U1��1��23�2@�U2M�2Z�2g�2t�U2��2��2��2��U2��2��2��2��2��2��33�����M�3Z�3g�3t�3���3��3��3��3���3��3��3��3���3��43�4@�4�M�4Z�4g�4t�4���4��4��4��4���4��4��4��4���4��53�5@�5�M�5Z�5g�5t�5���5��5��5��5���5��5��5��5���5��63�6@�6�M�6Z�6g�6t�6���6��6��6��6���6��6��6��6���6��73�7@�7�M�7Z�7g�7t�7���7��7��7��7���7��7��7��7���7�����Pv�U�B �@�09r�
�PV���A x� �0R���  ��BM�@RP�`�4Q_�PR�@[U�AR��D�SMC��E2F_�U��=A�QYSL|�P�@ �  � ֲ>g�������iD��VALU>e�pL��A�HFZAID_L����EHI�JIh�$FILE_ ��D�dc$Ǔ%`XCSA�Q� h�0!PE_BLCKz�.RI�7XD_CPUGY!�GY �Ic�O
T�Y.���R  � �PW`�p���QLA�n�S�Q�S�Q�TR?UN_FLG�U�T �Q�TJ��U�Q�T�Q�U�H��T`�T	 dw�T2L�_LIz��  �pG_�OT�P_ED�IU� 
/`�`7c� ?bة�pBQh��� ��TBC2 �! �%�>��P��a�7a�FTτ�d݃TDC"�PA�N`�`M�0�fL�a�gTH��U��d��3�gR�q�9�ER�VEЃt݃t	���a�p�` "Xw -$EqLENЃ0Rt݃Ep�pRAv��&Y@W_AtS1Eq�DM2�wMO?Q�S���pI�.B�A�y�4Ep��{DE�u��LACE �CCC�.B��_MA��v��w�GTCV�:��wT,� ;�Z�P���s�~��s*�J�A�M�����J���uā�uQq2ѐ���݁�s�JK��VK�������	���J����J�J�JJ�AAL��<��<�6��:�5�cm�N1a�m�,��
DL�p_\�Űѐ�a�CF
�# `�0G�ROU�@J�Բ��N�`C^�ȐREQUsIRrÀEBUu��Aq��$T�p2"���Bp薋a	��d$ y\?@qhAPPR��[CLB
$H`N;�'CLO}`K�S�e`���u]`BCI�% �3�M�`�l��_MG񱥠C �"P�����&���BRK��N�OLD����RTM!O6a�ޭ��J6`�P>��p��p��pZ�(�pc��p6+�7+�<���QAq�d&� �lr��������PATH���������qx�����%0A��S�CAub��<���INFDrUC�p�q�C�KUM�Y�psP�� ��A q/ʤ�/�E�/��PAYLOA�J{2L�0R_AN�ap�L�Pz�v�jɆ����R_F2LSHRt��LO{�R����|���ACRL_�q �����b��H�@B�$H��"�FLE�X>��aJ�f' P(��o�o+�p?q}JDu( :Q cv�p����f��po��|F1���-�@�����]�E� �*�<�N�`�r����� 4�Q�������A�c����ɏۏ���T��2�X :A�������� ��)�;�?�H�6�Z��c�u�������J��) ��`��˟ݟ�`�0cATF�𑢀EL��(a��J�(��J�E۠CTR��A�T�N�1�HAND_VBB>ѯ@�7* $��F2���d��CSW>�SATB���+� $$M �����0ˡ�ڡ������A�@g����AD)��A���@˪A٫AA� ��`P˪D٫�D�PȰG�P�)S�Tͧ�!ک�!N�DY�P9����#%��Fp ���Ѫ���i����������P3�<�E�N�W��`�i�r� =Ґe,1 ��ԓ� n�5<m��1ASYMص.@	�ض+A������_`��	���D� &�8�J�\�n�Ju�&���ʧC�I��S�_VI�o�Hm��@V_UANVb�@
S+��J� "RP5"R��&T��3TWV �͢���&��ߪU��a/�7Ԣ1�`HR`�ta-��QQ�1�DII��O�T���QN��. ; *"IAA*���$aG�2C2cJ��$��I��P / �� �ME��� Mb�R4AT�PPT@�@� ��ua����PАl@zh�a�iT�@��� $DUMMY}1E�$PS_D�RF��P$�fn3�FLA��YP����b}c$GLB_�T��Uuu`1�	�8��EQa0 X(����ST����SB}R�PM21_V��T$SV_ER��1O_@KscsCLpKreA��O'b�PGL�@;EW��1 4��aW$Y,Z,W�s怯��AN`©�q]U�u2 ��N�pސ@$GIU}$�q �p�s�p���3 L���v^B}$�F^BE�vNEARʖ�NK�F8���TAsNCK�w�JOG���� 4`$JOOINT�� $pސqMSET��5 E �wE�H�� S��
`�� ��6� � MU��?���L?OCK_FO�����PBGLVHGL��TEST_XM�>���EMPt���8�r̀$U�ГrF��22���s,�3��h�Ҁ,�1MqCE��|�sM� $KAR��}M�STPDRA�pj�a�VEC��{�e�kIU,�41�HEԀOTOOL㠓V�;RE��IS3����96N�A�ACH���E5��O�}c�d3����pSI.�  �@$RAIL_B�OXE��ppRO�BO��?�pqHOWWAR*���`�ROLM�bB����S��
�5���O_F�� !ppHTML	5�Q����Hb�pڑ��7m��R
��O��8���v�z���vOU��9 tpp(�14A�̀���PO֡%PIP��N��
�ڑS�,������CORDED0Ҁް̠5�XT��q�) �� O4` :o D pOBP! "Ҁ{�j��cpj�^@�$SYSj�ADR�#�Pu`TCH� o; ,��EN�R*Z�Aف_�t״�zbd�PVWVAPa?< � p��r��UPREV_RT~]1$EDIT�_VSHWR�7v(;���q�@D_`#�R�+$HEA�DoA�Pl�A$�K�E�q�`CPSPD���JMP��L�UMg�TR��d=r�TO�϶I�S#Ci�NE��$_TIC�K�AMXѭ ��H=N-q> @t������_GP��[�gSTYѲ�LOqPc��Ҩ�?�
�MGݵ%$���t=7pS !$Q��da��e!`�fP�0�SQ�Ud� ��b�ATER�Cy`,� S�@ �pCp����d�ė�%Oz`mcO�IZh�d�q�e�aPRM�0�a8����PUQH�g_DO=�ְXS���K�VAXIg�f�1�UR� ��$#��ȕ��� _����ET���Pۂ���5f�Fd�7g�A�!�1�d�9�2;"rSR|Al�о�� �#��5��#��#� )#�)i�>'i�N'i� ^&{����){����2��	C����C��WOiO{O܍D�qSSCp 7B hppDS(�k�f�`SP`�ATL ��I���¼bAD�DRES��B'�S�HIF��"�_2C�H#��I&p���TU&pI� C>��CUSTO����V��IbDȲ�,��0
�
_ED8U�R`E \����A�f�7��tC�#�	���F��irt�T�XSCREEl�Fz�P��TINA�s��p��t���Q_��0G T��fp,� ��eqBp&uᦲu�$#�RRO'0R���}��!Cd��0UE��H# ��0���`S�q��'RSM�k�UV����V~!�PS_�s�&C �!�)�'C��Cǂz"�� 2G�UE©4Ibvr�&8�GMTjPLDQ��Rp����R�BBL_�W��`R`J �f�>2O�qJ2LE�U3"��T4RIGH^3B�RDxt�CKGRĦ`�5TW��7�1WIDTH�H�Bb���a���T�UIu�E9Y��QaK d�p���A�J�
�4�BAC�KH��b�5|qX`F�OD�GLABS�?�(X`I�˂$UAR(�9@#p�0^`H4!� L 8�QR�_k��\B_`R�p͂�����HBO�R`M���w0Uj0�CRۂM�LUM�C��� GERV� �0P<�j�4NV`��GE=B0#���]�t�LP�E��	E��Z)Wj'Xz�'XԐ&Y5$[6$[7$[8	R���3�<��ԾfԑŁS��M��1USR�tO �<��^`U�r�rF�O
�rPRI��mx����PTRIP�m�UNDO��P�p��`m�4��l�,�#���� qQWB�P7�G s�aTf�H�RbOS�a�gfR��:">c��.qR`��s�~�b*� >c	UQ.qS�o�o�#R�)�>cOFF���pT� �cOp 1�R�t/tS�GU��P.q��JsETw�1�SUB*� f�E/_EXE��V��>c�WO>� U�`�^g��WA'��P�qz!@� V_DB�s��pEBSRT�`
�V0�Q�r��OR��u'RAU��tT�ͷr�q_���W |%��͸OWNA`޴$GSRCE � ��D��<\��MPFIA�p��ESPD������C���Gƒ�)�5��!GX `�`�r޴�n��COP�a$*�C`_w������rCT�3�q���qƒ ���@� Y"SHADOW�ઓ@�?_UNSCA��@���4M�DGDߑ��E�GAC�,��PP�G�Z (0N�O�@�D<�PE�Bf��VW씸�RG���![ � ��VqEE#��ڒANG�$���c薴cڒLIM_X�c��c� �����#��`� 퐾�VyF� �s�VCCj�j��\ՒC{�RAl�p����RpNFA�i�%�E��Z`�G� ^0[�C`DqEĒ��� STEQ1 ���@�ꁻ@I��`+0�����`����P_�A6�r���K��!]�� 1Ҡ��� ��\��сCPC�@]�GDRIܐ\�͑V#�耴��D�TMY_UBY�T���c��F!����Y��$���P�_V�y��LN�BMvQ1$��DEY��cEX�e��MU��5X�M� US�����P_R����P� ߖ=G��PACIr�ʐ f�ᔟ��c�´c���#B�EqB��aWrB�����^ ܀GBΐPK��)�D�R~`�`�_�0�@3!�1zr	4�e�R�SW��p��Yp��S�6�O�Q�1Ah� X�#�E�UE���Yp��C�HKJ�`�@p���U� �EAN�ٖp�pX���MRCV�!a ���@O��M�pCL	p��s����REF*7 
��������/��P�ڀ@���@��b��֗�_ Y��ژ��ۣ��Q$3ಲ���?��$b �����%���Q��$GROU� �c���d��ʠ]��I2^00��U` 0_�IX,�o � ULա`���C&�rAaB�?�NT����$����A���Q��K�L����õ��A����Q��T a$c �t�`MD�p8�HUح��SA��CM�PE F  _��Rr�p@����X�S	qVGF/�b#d/, &�@M�P^0۰UF_C !���z �ROh0"+���@8���0C�UREB�f��RI��
IN�p �����d��d��ca�INE�H�y��0�V�a-�걗�3�W �������C��i�LO�}�z�@0�!�QNSI��݁���c�$&�c$&.�X_PE:-YW+Z_M�ڒ�W�I�$�" �+R܃'rRSLre I�/�M
`�R
E�C7�Gd�۰�̵� ��q����u��Ȑ ������S_P�VnP� ��IA�vf ]�~pHDR�p�p�JO�P��$�Z_UP��a_�LOW�5�1J�dAn��LINubEP?�@tc_i�1�1���@�G�1@d�0W�xg{ 5X�PATHP= X�CACH$��]E��yI�A��{�C�)�ID3FA�ETD��H��$HO�pղb@�{�d6�F����<��p�PAGE�䁀�VP�°�(R_SI	Z��2TZ3�-X�0U̲q�MPRZ��IM5G���AD�Y��MRE��R7WGP���8�p��ASYN�BUF�VRTD��U�T7Q�LE_2�D-��U��`CҡU�1��Qu��UECCU��VEM��]EDb�GVIRC�Q�U�S��B�Q�LA��p�N�FOUN_�DIAuG�YRE�XYZ�cE�WѴh8�dpq2a`T��2�IM�a�V�|be��EGRABBr��Y�a�LERj��C4���FC-A�65a04x��7u$� BE���h��`�CKL�AS_@l�BA��N@i�  G��T��� @�ݲմ$BAƠwj A�!q�eb��uTYS p�H����2��I�t:bt�f��B)�EVE�����PK���fx��GI�pNO��2����q�HO����k � ����
8�Pi�S��0ޗ��RO��AC�CEL?0=���VR_�U7@�`��2�p�6�AR��PA��̎�K�D��REM_B6ut N�JMX ��l�t�$SSC��U �
�#���QN@m� � �S�P�N�S���LEX�vn =T�ENAB 2¼W@��FLDRߨF�I�P�t�ߨ(Ğ��� �VP2HFo'� ��V
Q MV_PI��8T @󐉰�F@�Z�+�#��8�8�#��GAB���LO9O��JCBx��w�"SCON(P�PLCANۀ�Dp�3F�d�v�9PէM��Q ;����SM0E�ɥ�8�ɥWb72$`<�8T̸�,`RKh"ǁVAsNC���1R_Ou N@p (�-#<#c���c2A04w�A/�N@q 4�������`	�^�o�r h�n���1^�&OFF�`|�p�`��`�DEeA�
�P,`SK�D�MP6VIE��2q� w��@���rs �< {���4��h�r{7��D���
ѯCUST�U��wt $G�TIT1�$PR\��O�PTap ��VSF�йsu�p�0`r&��̑SMOwv�I�|�ĄJ������eQ_WB��wI����� @O3�@�XVR�xxmr��T����ZABC���y op����)�
�� 
�ZD$�CwSCH��z Lu� ���`�2�%PC ��7PGN ��<��A��O_FUNH��@�̐7ZIPw{I��KLV,SL��~�)P��ZMPCF��|���E����X�DMY'_LNH�=�4D�� ~��} $�A�� ]�CMCM� C�,SC&!��P�� �$J���D Q�������������a_�Q,2����UX�a>\�UXEUL��a ������(�:�(�J���FTFL��w�7	�Z�~Zp+ڦ6� �p��Y@D�p  8 �$R�PU��> EI3GH����?(�i���M���et� �0a�����$B�0�0�@�	�_SHIF,D3-�RVV`F�@��	$5��C�0��&! ������b
�sx��uD�TR��V�̱SPH���!�C ,��������4A��RYP��%������%�ː"�%!W  �H�(UN0���"�2������ɒ�q0G�SPDak�� ��P��O����0X��Ѱ�"!�NGVER`q �iw+I_�AIRPURGE�  i  �i/�F`E�Tb� ��+1h2ISOLC�  �,�"ːDː�!�%��P+�_/�*OB��Dm�?�@�!H771  34n?�?@�9� `�E/#�)x� �S232�� 1�i� LT�Ek@ PENDA`�341 1D3<�*? Ma�intenanc�e Cons B��? F"O,DNo UseMJOOnO��O�O�O�O2�2NPQO;/" 19%�1;CH=� �.ː�		9Q_!U�D1:___RSM�AVAIL/�/%��A!SR  ��+��H�_�P1�TVAL.&���P(.r�YVL�}� 2i��� D��P 	�/_oUQNo�orc i�o�g�o�o�o�o�o *,>tb� �������� :�(�^�L���p����� ��܏ʏ ��$��H� 6�X�~�l�����Ɵ�� �؟�����D�2�h� V���z��������ԯ 
���.��R�@�b�d� v�����п��������(�N�<�r�i�$�SAF_DO_PULS. jQp��F��CA� �/%�&�0SCR �`X�_�0�0�
	14�1IAIE���b vo$�6�H�Z�l� ~�ߢߴ���������V�HS��2%�$��0�d%�@�rb��� @�"k�}��ȡ�T�h� J`��_�_ @��T7 ������#�0�T D��0�Y�k�}��� ������������ 1CUgy�O�Ef������  �5;�o��� 1p�U�
�?t��Di��������
  � � �*������gy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�?@�?OO%O7O<A��� `OrO�O�O�O�O�O�O �O?O�_._@_R_d_ v_�_�_�_�_�Q _�R0MJTo!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏJO� �'�9�K�]�o����� ��_ɟ۟����#� 5�G�Y��_�U�_�ҙ� ����ϯ����)� ;�M�_�m��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f�;�?�q߮����� ������,�>�P�b�t���������p��������Y���	123�456781h!B!����
F��������� �������� �� ;M_q���� ���%7I [l*����� ��//1/C/U/g/ y/�/�/�/n��/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?O�/ )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_O_�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�op_�o�o �o/ASew �������� �o+�=�O�a�s����� ����͏ߏ���'� 9�K�]���������� ɟ۟����#�5�G��Y�k�}���������s�կ�w���0��L�CH  Bp�w�   �=�2��� }� =�
���  	�o�ί��ǿٿ$���r������@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖ�%Ϻ������� ��&�8�J�\�n�� ��������������"�Q�*�����;�<�M���D���  �]�w�*�Z�>��t  d������*�`*��$SC�R_GRP 1�*P3� �� �*�� 6�	 /�
 ��<�+*�'UC�|@��y�yD� W�!�y��	M-10iA�/7L 1234�567890��v� 8��MT� �� �
�	L��,	Č� N
�@��Y���y�
M_	P������ ,��H�
 ���1/@A/ g/y/H�ߙ!T/�/�P/�/3��+���/B��S��,?*2C4&Ad�R?  @s�j5N?�7?��7&2R��?}:�&F@ F�` �2�?�/�?�?OO-O SO>OwObO�O=j1�2`�O�O�O�O�DB��O �O;_&___J_�_n_�_ �_�_�_�_o�_%o�@5j�eSgxo6����uo�o�b�1�B�8K`�oh0�4j9j9B� w�$Y̯@HtCA�Nhcu�/�%pp�drsq �����z�q�x� �� (&�*�2�D�V��oz�e�������EC�LVL  �����iqpQ@��L�_DEFAULT� ���s�փHOTST�R�qq��MIPO/WERF��H��WFDO�� �RVENT� 1ɁɁ� �L!DUM_E�IP�����j!?AF_INE‧����!FT}�֞䝟��!-/� ���F�!RPC_OMAING�)��5����Y�VISb�t�����ޯ!TPѠP�Uկ��dͯ*�!
�PMON_PROXY+���e�v���D���fe�¿!R?DM_SRVÿ��9g���!R,*ϲ��h��Z�!
[�M䍿��iIϦ�!R�LSYNC�����8����!ROS�|���4��>�!
�CE�MTCOMd?ߓ�k-ߊ�!	S�OCONS�ߒ�ly����!S�WASR�Cݿ��m��"�!NS�USB#n�>n�!STMC�����o]�����ѳ������,���P�V�ICE_KL ?%d�� (%SVC�PRG1S�����2�������3������4�������5��6;@��7ch��$���9����%� �������0�� ��X�����-� ��U���}���  /���H/���p/�� �/��F�/��n�/ ��?��8?��� `?��/�?��6/�?�� ^/�?��/X�j��q� ��#OhO��lO�O{O�O �O�O�O�O�O _2__ V_A_z_e_�_�_�_�_ �_�_�_oo@o+odo Oo�o�o�o�o�o�o�o �o*<`K� o������� &��J�5�n�Y���}�एȏ���^�_DE�V d���MC:�4��~�GRP 2d��
@�bx 	_� 
 ,V�I� �s�Z��������� ���ߟ��@�'�9� v�]�������Я���� ۫Y��.��R�9�v� ��o�����п_�ǿ� �(��!�^�Eς�i� �ϸ��a��ϥ���� 6��Z�l�Sߐ�wߴ� �߭������ ��D� +�h�O����U����� ���������R�9� v�]������������� �������^� i�����  �)>�bI�� ����I/� :/L/��p/W/�/{/�/ �/�/�/�/?$??H? /?l?~?e?�?��?�? �?�?�? O2OOVO=O zO�OsO�O�O�O�O�O 
_�O.__R_d_�?�_ k_�_�_�_�_�_oo �_<o#o`oroYo�o}o �o�o�o�o�o�o}_ Jn�g��� ����"�	�F�X� ?�|�c�������֏��d �X�ZI6� r 	 @�Z��0�+A�����dBjBA�=��������B����AZ.�AĊ��+�A.��Q�B����5�\��i6�A��u��'����%�Ꮛ�%P�EGA_BARR�A_ESTEIR�A������� ʑ&�ʕڟ�ҟ���0,��P�^�%�����  >�`�:���ޯ̯ ��&�h�M������ n�������ڿȿ��@� %�d��X�F�|�jό� �Ϡ������<���0� �T�B�x�f߈���� ��߮����,��P� >�t�ߛ���d���`� �����(��L���s� ��<�����������  ��$f�K��~l ������># b�VDzh�� ������/ R/@/v/d/�/��/ / �/�/�/???N?<? r?�/�?�/b?�?�?�? �? OOOJO�?qO�? :O�O�O�O�O�O�O�O ROxOI_�O"_|_j_�_ �_�_�_�_*_oN_�_ Bo�_Roxofo�o�o�o o�o&o�o>, Ntb��o��o� ����:�(�J�p� ����`�ʏ���܏ � �6�x�]�o�&�H� "���Ɵ���؟�P� 5�t���h�V�x�z��� ¯���(��L�֯@� .�d�R�t�v����� � �$�����<�*�`� N�p�ƿ쿽������� ����8�&�\ߞσ� ��L߶�H�������� ��4�v�[��$��|� ����������N�3� r���f�T���x����� ����&�J���>, bP�t����� ���:(^L ����r��� � /6/$/Z/��/� J/�/�/�/�/�/�/�/ 2?t/Y?�/"?�?z?�? �?�?�?�?:?`?1Op? 
OdORO�OvO�O�O�O O�O6O�O*_�O:_`_ N_�_r_�_�O�__�_ o�_&oo6o\oJo�o �_�o�_po�o�o�o�o "2X�o�oH �������` E�W��0�
�x����� ҏ����8��\��P� >�`�b�t�����Ο� ��4���(��L�:�\� ^�p����ͯ��� � �$��H�6�X���ԯ ���~�ؿƿ��� � �Dφ�kϪ�4Ϟ�0� �����������^�C� ���v�dߚ߈ߪ��� ����6��Z���N�<� r�`��������� 2��&��J�8�n�\� �����������~��� "F4j����� Z����� B�i�2��� ����/\A/� 
/t/b/�/�/�/�/�/ "/H/?X/�/L?:?p? ^?�?�?�?�/�??�? O�?"OHO6OlOZO�O �?�O�?�O�O�O_�O _D_2_h_�O�_�OX_ �_�_�_�_
o�_o@o �_go�_0o�o�o�o�o �o�oHo-?�o �o`�����  �D�8�&�H�J�\� �������ݏ���� ��4�"�D�F�X���Џ ���~��֟���0� �@�������̟f��� ���ү���,�n�S� ������������� ο�F�+�j���^�L� ��pϒϸϦ����� B���6�$�Z�H�~�l� �ߴ�����ߤ���� 2� �V�D�z�ߡ�� j��f���
���.�� R���y���B������� ������*l�Q�� �r����� D)h�\J� n���
0/@ �4/"/X/F/|/j/�/ ��//�/�/�/
?0? ?T?B?x?�/�?�/h? �?�?�?�?O,OOPO �?wO�?@O�O�O�O�O �O�O_(_jOO_�O_ �_p_�_�_�_�_�_0_ o'o�_ o�_Ho~olo �o�o�oo�o,o�o  02Dzh��o �����
�,� .�@�v�����f�Џ ������(�~��� u���N�����̟��� ޟ�V�;�z��n� � ~�����ȯ���.�� R�ܯF�4�j�X�z��� ��Ŀ��*����� B�0�f�T�vϜ�޿�� ό�������>�,� bߤωߛ�R�t�N߼� ������:�|�a�� *���������� �T�9�x��l�Z��� ~���������,�P� ��D2hV�z� ���(�
@ .dR����x �t�//</*/`/ ��/�P/�/�/�/�/ �/??8?z/_?�/(? �?�?�?�?�?�?�?O R?7Ov? OjOXO�O|O �O�O�OO�O_�O�O �O0_f_T_�_x_�_�O �__�_o�_oo,o boPo�o�_�o�_vo�o �o�o(^�o ��oN���� � ��f�]��6��� ~�����؏Ə��>�#� b��V��f���z��� ��ԟ���:�ğ.�� R�@�b���v����ӯ ������*��N�<��^���Ư������$SERV_MA_IL  �����ʴOUTPU}Tո�}@ʴRV 2j�>ǰ�  (r�������=�ʴSA�VE���TOP1�0 2� d? 6 rƱ�� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b�0t�����n�YPY���FZN_CFG ;j��=���J���GRP 2���g� ,B �  A �D;�� B �  B�4=�RB21�I�HELL�� j�e�)�*�=����>�%RSR�� ����&J 5G�k�������.�  ���/>/P/"\/ ��X/z"{ �U'&"2�dh,g-�"�EHK 1S �/�/�/�/#?L? G?Y?k?�?�?�?�?�? �?�?�?$OO1OCO??OMM S�O�DFTOV_EN�BմƱe��"OW_?REG_UI�O��IMIOFWDL�~@�N�BWAIT�B�)��V��F��YTIM�E��G_VA԰_�A_UNIT�C~VeɻLC�@TRY�G�e�ʰMON_ALIAS ?e�I%�he��oo&o 8oFj�_io{o�o�oJo �o�o�o�o�o/A Sew"���� ����+�=��N� s�������T�͏ߏ� ����9�K�]�o��� ,�����ɟ۟ퟘ�� #�5�G��k�}����� ��^�ׯ�����ʯ C�U�g�y���6����� ӿ忐����-�?�Q� ��uχϙϫϽ�h��� ����)���M�_�q� �ߕ�@߹������ߚ� �%�7�I�[���� �����r������!� 3���W�i�{���8��� ����������/A Se����� |�+=�a s��B���� /�'/9/K/]/o// �/�/�/�/�/�/�/? #?5?�/F?k?}?�?�? L?�?�?�?�?O�?1O COUOgOyO$O�O�O�O �O�O�O	__-_?_�O c_u_�_�_�_V_�_�_��_ooc�$SM�ON_DEFPR�OG &����Aa &�*SYSTEM�*obg $J�O0dRECALL� ?}Ai ( ��}tpdis�c 0=>10.�109.3.13�2:21064 �4 �l�e0�`87�40bo�o�o	w}�tpconn 0 �o�o�o[mw�8copy fr�s:orderf�il.dat v�irt:\tmpback\�o7pV���}/�rmdb:*.*���^��p���t3x�t:\ &���8�7pQ����
p4��a����Kvӏ�d�v���}?�:p�ickup_ba�rra_este�ira.tp)�emp7�6qܟ� �v�=����torno@��˟۟l�~�x6�lace1�C�P�U�����~<�sumir+���њۯl�~�������prens ��G�Z������+� ��ؿi�{�� �;�D� V����ό���1�G��� e�w�
��-�?�R��� ����,ϵ���a�s� ���3��N������ ߩ߻�L�]�o����߀%�7��߉�����w
�xyzrate 11 ������]o4�u61=7p <N���� �]o�������0y V����.y�� _/q/�/@/:/L/�/ �/?/&/�/�/	?m? ?�/�/6?H?Z?�?�? ?"?�?�?�?iO{O�? �?2ODOVO�O�OOO �O*_�Oe_w_
_�.� >_R�_�_o��_�� �_aoso�o�+8oN� �o�o���o�oL] o��_�_/o�_�� �o$o�Ho�k�}� �o�o5�oX����  ��D֏g�y��� �>�T����������@�ҟc�u��� �$�SNPX_ASG 2�������  �0��%���Я  �?���PARAM� ���� W�	��PӤ��9Ө$�������OFT_KB_CFG  ӣ�����OPIN_SIMW  ���}����������RVNO�RDY_DO  �)�U���QST_P_DSBi��|ϐ�SR �� � &#�D�O��O�:�TOP_ON_ERRʿ��o��PTN ��ޢ��A��RI?NG_PRMy�ܲ�VCNT_GP �2��!���x 	���ϗ���#��G����VD��RP 1	��"�8Ѩ�*߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�}�z��������� ������
C@R dv������ 	*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?[?X?j?|?�?�?�? �?�?�?�?!OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLosopo�o �o�o�o�o�o�o  96HZl~�� ������ �2��D�V�`�PRG_CoOUNTJ���N{�ENB��}�M���L���_UPD 1}'�T  
k� �����"�K�F�X�j� ��������۟֟��� #��0�B�k�f�x��� ������ү������ C�>�P�b��������� ӿο����(�:� c�^�pςϫϦϸ��� ���� ��;�6�H�Z� ��~ߐߢ��������� �� �2�[�V�h�z� ������������
� 3�.�@�R�{�v����� ��������* SN`r���t��_INFO 1��Ҁ� 	� ��3@�ub?���?#Ҹ�D�v:� B��L���A��BA�V������>>@ A�� ?�| @�| ?M @��9 ¶���C�y�C��K��3���?��B� ����YSDEBUG������ dՉ�S�P_PASS���B?+LOG u���  � 99�  �с�UD1:\;$<�<"_MPCA-�H�/�/�x!�/ �~�&SAV D)`��%d!|"�%�(�SV�+TEM_T�IME 1D'��� 0Ҁ<΄��(�/�3Q3MEM�BK  �с�d d/�?�?�<X�|Ҁ� @�?C��O:OJLOmOzI,�J
! %@p1�O �O�O�O"3 __$_6_H_Z_l_ �n_�_�_ �_�_�_�_�_o"o\�e1oVohozo�o�o�o �o�o�o�o
.@�Rdv���O5SK�0�8���?���VF=� "�H2OJ�AJ� l�\C�Ah\O����(�O!��O�я�����O!�� �!�j�TO^�p���v_��U����ӟ���	��� $�C�7og�y� ��������ӯ���	� �-�?�Q�c�u�����������T1SVG�UNSPD%% '�%��2MOD�E_LIM �a9"ܴ2�	� �D-۵ASK_OP�TION �9!�F�_DI ENB�  U�%f�BC�2_GRP 2!@�u#o2��N��C�����ԼBCCFG 3#��*< #6���`�@I�4�Y� �jߣߎ��߲����� ����E�0�i�T�� x������������ /��S�>�w����6u� ��u�����c���	 B-f�.��4[ � ������  02Dzh��� ����/
/@/./ d/R/�/v/�/�/�/�/ �(���/?&?8?J?�/ n?\?~?�?�?�?�?�? �?O�?4O"OXOFOhO jO|O�O�O�O�O�O�O __._T_B_x_f_�_ �_�_�_�_�_�_oo >o�/Voho�o�o�o(o �o�o�o�o(:L p^����� ��� �6�$�Z�H� ~�l�������؏Ə�� � ��0�2�D�z�h� ��To��ȟ���
��� .��>�d�R������� z�Я�������(� *�<�r�`��������� ޿̿���8�&�\� Jπ�nϐϒϤ����� �ϴ��(�F�X�j��� ��|ߞ��߲������ ��0��T�B�x�f�� ������������� >�,�N�t�b������� ����������:( ^�v����H ���$HZl :�~����� ��2/ /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?P?R?d?�?�? �?t�?�?OO*O�? NO<O^O�OrO�O�O�O �O�O�O__8_&_H_ J_\_�_�_�_�_�_�_ �_�_o4o"oXoFo|o jo�o�o�o�o�o�o�o �?6Hfx� �������v&���$TBCSG_�GRP 2$�u��  ��&� 
 ?�  Q�c�M���q���������ˏ��*�1�&~8�d, �F��?&�	 HCA������b��CS�B�I������V�>��ͪ�n��쌟ԝB��333,��Blt�����r�AÐ�fff:�L�.�C����l�?����G�w�R���A&��̧�����@��I��-���
�X��u�@�R�����̻������	V3.00>I�	mt7����*� �%��ֶY�_�@ff&� &��H�� N� �O� ; ����� ϏϬ��*�J21�'8���Ϥ�CFG )��uB� E�������d���#��#�I�W��pW�}� hߡߌ��߰������ ��
�C�.�g�R��v� ��������	���-� �Q�<�u�`�r����� ������I�cp" 4��gRw��� ���	-?� cN�r��&�� ����/</*/`/ N/�/r/�/�/�/�/�/ ?�/&??J?8?Z?\? n?�?�?�?�?�?�?O �? OFO4OjOXO�O�O `�O�OtO�O_�O0_ _T_B_x_f_�_�_�_ �_�_�_�_�_,ooPo boto�o@o�o�o�o�o �o�o�o(L:p ^������� � �6�$�F�H�Z��� ~�����؏Ə���� 2��OJ�\�n������ ��������
�@� R�d�v�4��������� ί����ү(�N�<� r�`���������ʿ̿ ޿��8�&�\�Jπ� nϐ϶Ϥ��������� "��2�4�F�|�jߠ� �����߀��� �߼� B�0�f�T��x��� ����������>�,� b�P���������v��� ����:(^L �p�����  �$H6lZ| ������/� / /2/h/�߀/�/�/ N/�/�/�/
?�/.?? R?@?v?�?�?�?j?�? �?�?�?O*O<ONOO O�OrO�O�O�O�O�O �O _&__J_8_n_\_ �_�_�_�_�_�_�_o �_4o"oXoFoho�o|o �o�o�o�o�o�/$ 6�/�oxf��� �����,�>�� �t�b�������Ώ�� 򏬏��&�(�:�p� ^���������ܟʟ� � �6�$�Z�H�~�l� ������دƯ��� � �D�2�T�z�h��� Jȿڿ������
�@� .�d�Rψ�vϬϾ��� �Ϡ������*�`� r߄ߖ�Pߺߨ����� �����&�\�J�� n������������ "��F�4�j�X�z�|� ������������0 B�Zl~(�� �����,P bt�D�������   #� &0/"�$T�BJOP_GRP� 2*��  ?�&i	H"O#,V,��w�� �� �=k%  Ȫ �� �� �$ �@ g"	 �CA���&��SC���_%g!�"G���"k��/�+=��CS�?ϙ�?�&0%0CR  B4�'??J7�/^�/?333�2Y&0<}?�:;��v 2�1)�0-1*20�6?�?�20��7C�  D��!�,� BL���OK:�Z�Bl�  @pB@�� s�33C�1 �?gO ' A�zG�2jG�&�)A)E�O�J;��>|A?�ff@U@�1�C�Z0zjO�Oz@����U�O�$fffx0R)_;^;xCsQ?ٶ4)@�O�_tF�X�_J\EU�_�V:�t	-�Q(B�*@�Ooh �&-h$oZGLo6oDoro �o~o8o�o�o�o�o 3�oRlVd���V4�&`�q�%	�V3.00m#'mt7A@�s*�l$�!�'� E���qE���E��]\E�HF�P=F�{F*�HfF@D�FW��3Fp?F��MF���F��MF��F��şF��F��=F���G��G.8�C�W�RD3l)D���E"��E�x�
E��E��,)FdRF�BFHFn� F���F��MF��ɽF�,
G�lGg!G�)�G=��G�S5�GiĈ;��
;�o�|U& : @Xz&/T��&"�?�0��&=;-ESTPARS  (a E#�HRw�ABLE ;1-V) @�#�R�7� � �R�BR�R�'#!R�	R�E
R�R���!R��R�R���RD	I��`!��ԟ���
�r�Oz����������̯ޮ��Sx�^#  <�����ÿտ���� �/�A�S�e�wωϛ� �Ͽ�������;-w�{� _"��6��1�C�U����%�7�I�[����N�UM  �*`!� $  ��m����_CFG .����!@H IMEBF_TT}���^#��G�VE10m�H�]�G�R 1/��' 8�" �� �A�  ����� ������� �2�D�V� h�z������������� /
e@Rhv ������� *<N`r�� ����'///]/ 8/J/`/n/�/�/�/�/�r���_��t�@~��t�MI_CHAN�S� ~� !3DBGLVLS�~�s�$0�ETHERAD �?��w0�"���/�/�?�?l�$0RO�UTq�!�!��4�?�<SNMAS�Kl8~�}1255.2E�s0OBOTO�st��OOLOFS_D�I}��%V9ORQCTRL 0���#��MT�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo&l�O�Io8omoq�PE_D�ETAIJ8�JPG�L_CONFIG� 6�ᄀ�/cell/$C�ID$/grp1�qo�o�o/壀 �?Zl~���C ���� �2��V� h�z�������?�Q�� ��
��.�@�Ϗd�v� ��������M����� �*�<�˟ݟr���������̯@�}a��� &�8�J�\���^o��c��`���˿ݿ��� Z�7�I�[�m�ϑ� � �����������!߰� E�W�i�{ߍߟ�.��� ���������A�S� e�w����<����� ����+���O�a�s� ������8������� '9��]o�� ��F���# 5�Yk}������`�User View �i�}}1234567890�//,/�>/P/X$� �cx/���2�U�/�/�/�/ ??s/�/�3�/b? t?�?�?�?�??�?�.4Q?O(O:OLO^OpO�?�O�.5O�O�O�O@ __$_�OE_�.6�O ~_�_�_�_�_�_7_�_�.7m_2oDoVohozo�o�_�o�.8!o�o�o�
.@�oagr �lCamera��o����� �ޢE�*�<� N��h�z��������I  �v�)��$� 6�H�Z�l�������� ��؟���� �2�Y��vP9ɟ~������� Ưد���� �k�D� V�h�z�����E�W�I 5����� �2�D�� h�zό�׿�������� ��
߱�W�ދ��X�j� |ߎߠ߲�Y������� E��0�B�T�f�x�� �ulY���������
� ���@�R�d������ ����������W� iy� .@Rdv�/�� ���*< N��W��i���� ����/*/</� `/r/�/�/�/�/as9F/�/??1?C?U? �f?�?�?D/�?�?�?��?	OO-O�j	�u0 �?hOzO�O�O�O�Oi? �O�O
_�?._@_R_d_ v_�_/OAO�p�{,_�_ �_oo)o;o�O_oqo �o�_�o�o�o�o�o �_�u���oM_q� ��No���:� %�7�I�[�m�NEa� ���ˏݏ���� 7�I�[���������� ǟٟ����ͻp�%�7� I�[�m��&�����ǯ �����!�3�E�� ��9�ܯ������ǿٿ 뿒��!�3�~�W�i� {ύϟϱ�X�����H� ���!�3�E�W���{� �ߟ������������<���  ��L� ^�p���������x�� ��   "� *�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/��  
��(  ��@�( 	  �/�/�/�/�/? ?6? $?F?H?Z?�?~?�?�?t�?�*2� �l� O/OAO��eOwO�O�O �O�O��O�O�O_TO 1_C_U_g_y_�_�O�_ �_�__�_	oo-o?o Qo�_uo�o�o�_�o�o �o�o^opoM_ q�o������ 6�%�7�~[�m�� �������ُ���D� !�3�E�W�i�{�ԏ ��ß՟�����/� A�S���w�����⟿� ѯ�����`�=�O� a�����������Ϳ߿ &�8��'�9π�]�o� �ϓϥϷ��������� F�#�5�G�Y�k�}��� �߳���������� 1�C�ߜ�y����� ��������	��b�?� Q�c������������ ��(�)p�M_�q������0@ A�������� ��#frh:�\tpgl\ro�bots\m10�ia4_7l.xml�Xj|��������.�� /1/C/U/g/y/�/�/ �/�/�/�/�//?-? ??Q?c?u?�?�?�?�? �?�?�?
?O)O;OMO _OqO�O�O�O�O�O�O �OO _%_7_I_[_m_ _�_�_�_�_�_�__ �_!o3oEoWoio{o�o �o�o�o�o�o�_�o /ASew��� ����o��+�=� O�a�s���������͏�ߏ�I |�<<  ?��4��,�N� |�b�������ʟ�Ο ���0��8�f�L�~�@��������������(�$TPGL_�OUTPUT �9����� $�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}ϏϡϠ������$����2�345678901��� �2�D�V�^� ���υߗߩ߻����� w����'�9�K�]���}g��������o� ����1�C�U�g��� u�����������}��� -?Qc��� ������) ;M_q	�� �����%/7/I/ [/m///�/�/�/�/ �/�/�/?3?E?W?i? {??%?�?�?�?�?�? O�?OAOSOeOwO�O !O�O�O�O�O�O_�O~� $$Ӣ ��OW=_o_a_�_�_�_ �_�_�_�_�_#ooGo 9oko]o�o�o�o�o�o �o�o�oC5g}���������}@��"�� ( 	 iW�E� {�i�����Ï��ӏՏ ���A�/�e�S��� w��������џ��� +��;�=�O���s�����Ƹ  <<\ޯ�)�ͯ�)� �M�_���ʯ����<� ��ؿ��Ŀ� �~�$� V��BόϞ�x����� 2ϼ�
ߤ���@�R�,� v߈���p߾���j��� ����<�߬�r�� ��������`� &�8���$�n�H�Z��� �����������"4 Xj��R��L ����|T f ��v��0 B//�&/P/*/</ �/�/��/�/h/�/? ?�/:?L?�/4?�?? n?�?�?�?�? O^?�? 6OHO�?lO~OXO�O�O O$O�O�O�O_2__ _h_z_�O�_�_J_�_��_�_�_o.o��)�WGL1.XML��cm�$TPOF?F_LIM Š�p����qfNw_SVy`  �t��jP_MON �:���d�p��p2miSTRTC�HK ;���f�~tbVTCOMP�AT�h*q�fVWV_AR <�mMx.�d  e�p��bua_DEFPROG %�i�%COLOC�A_BARRA_TORNO A|~�sISPLAY�`��n�rINST_M�SK  �| ~�zINUSER ��tLCK)��{QU?ICKMENM��toSCREl���~+rtpsc�t�)������b��_��S�Tz�iRACE_�CFG =�i�Mt�`	nt
?�~�HNL 2>�z���T{ zr@�R�d��v���������К�I�TEM 2?,�� �%$1234?567890�%�  =<�C�U�]��  !c�k�wp '���ns�ѯ5���� k������j�ů��� ����A�1�C�U�o�y� 󿝿I�oρ�忥�	� �-ϧ�Q���#�5ߙ� A߽�����e߳���� ��M���q߃�L��g� �ߋ����%�w� � [���+�Q�c���o� �������3��� {�;������G_�� ��/�Se.� I�m�� �=�a/3/�� ����k//�/�/ �/]/?�/�/�/?�/ u?�?�??�?5?G?Y? �?+O�?OOaO�?mO�? �?�OO�OCO__yO +_�O�Ox_�O�_�O�_ �_�_?_�_c_u_�_o �_Wo}o�o�_�oo)o ;o�o�oqo1C�oO �o�o��%��@[��Z��S��@��_��  �ے_� ����y
� Ï�Џ����UD1:\����q�R_GRP 1�A �� 	 @�pe�w�a���������ߟ͞�����ّ�>�)�b�M�?�  }���y�����ӯ ������	��Q�?� u�c���������Ϳ��	-���o�SC�B 2B{�  h�e�wωϛϭϿ��������e�UTORIAL C{��@��j�V_CONFIG D{����������O�OUTPUT� E{�����������%�7�I� [�m�������� ������%�7�I�[� m�������������� ��!3EWi{ �������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/��/??'?9?K? ]?o?�?�?�?�?�?�/ �?�?O#O5OGOYOkO }O�O�O�O�O�O�?�O __1_C_U_g_y_�_ �_�_�_�_�O�_	oo -o?oQocouo�o�o�o �o�o�_�o); M_q����� �yߋ����-�?�Q� c�u���������Ϗ� ��o�)�;�M�_�q� ��������˟ݟ� � �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i�{������� ÿտ���
��/�A� S�e�wωϛϭϿ��� ������+�=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� �����������1 CUgy���� ���	-?Q cu��������/�x��� $/6/ !/a/��/�/ �/�/�/�/�/??'? 9?K?]?�?�?�?�? �?�?�?�?O#O5OGO YOkO|?�O�O�O�O�O �O�O__1_C_U_g_ xO�_�_�_�_�_�_�_ 	oo-o?oQocot_�o �o�o�o�o�o�o );M_q�o�� ������%�7� I�[�m�~������Ǐ ُ����!�3�E�W� i�z�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'��9�K�]�o�~��$T�X_SCREEN� 1F8%  �}�~���������
����m&�� \�n߀ߒߤ߶�-�?� �����"�4�F��j� �ߎ���������_� ���0�B�T�f�x��� ���������� ��>��bt��� �3�W(: L^������ ��e/�6/H/Z/�l/~/�//�/�$U�ALRM_MSG� ?�����  �/���/�/)??M?@? q?d?v?�?�?�?�?�?��?O�%SEV  ��-EF�"EC�FG H����  ��@� � AuA   B���
 O���ŨO �O�O�O�O__&_8_�J_\_jWQAGRP �2I[K 0��	� �O�_� I_B�BL_NOTE �J[JT�G�l������g@~�RDEFPRO� �%�+ (%M�AIN _PLACE�W2n%OVoAo zoeo�o�o�o�o�o�o��o@�[FKE�YDATA 1K<�ɞPp jG���_������z�,(�����OI�NT  ]'�)�?DIRECT}@o��*�INg����[?CHOICEB���?[LISTƏ��8�RE INFO ��C�U�<�y�`��� ����ӟ����	��-���Q�c� ���/frh/gui�/whiteho?me.pngd���p��Ưدꯀ  |�point���0��B�T�f���{�direc������οl��{�in����0�B�T�f�q�{�choic��ϰ�����������{�lis��2�D�V�h�z�>��arwrgϲ� �������߉��)�;� M�_�q������� �������%�7�I�[� m������������� ����3EWi{ ������ �/ASew�� r������/!/ (E/W/i/{/�/�/./ �/�/�/�/??�//? S?e?w?�?�?�?<?�? �?�?OO+O�?OOaO sO�O�O�O8O�O�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5o�_Goko}o�o�o �o�oTo�o�o1 C�ogy���� P��	��-�?�Q� �u���������Ϗj�-܋�u�܏�@(�s��Q�c�r�,I����A�POINT�  ]��9� IR�ECTß�}�ND�؟�F�CHOIC�E���TOUCHUPG�H�s���~� ����߯�د���9� K�2�o�V�������ɿ���whitehom����%�7��I�X��poin��ߍϟϱ����ψ�i?/direc|���$�6�H�Z���/in �ϓߥ߷�����j���choic���� �2�D�V�h�k��t?ouchup�ߠ�������g��arwrg��"�4�F� X�j�a����������� ��w�0BTf x������ �,>Pbt ������/� (/:/L/^/p/�//�/ �/�/�/�/ ?׿�/6? H?Z?l?~?�?�/�?�? �?�?�?O�?2ODOVO hOzO�O�O-O�O�O�O �O
__�O@_R_d_v_ �_�_)_�_�_�_�_o o*o�_No`oro�o�o �o7o�o�o�o& �oJ\n���� E����"�4�� X�j�|�������A�֏ �����0�B�яf� x���������O�������,�>�ټL�}�����u�@����q���ͯ��,�� ����"�	�F�X�?�|� c�������ֿ����� �0��T�f�Mϊ�q� �ϕ����������,� >�?b�t߆ߘߪ߼� ˟������(�:�L� ��p�������Y� �� ��$�6�H���l� ~�����������g���  2DV��z� ����c�
 .@Rd���� ���q//*/</ N/`/��/�/�/�/�/ �/�//?&?8?J?\? n?�/�?�?�?�?�?�? {?O"O4OFOXOjO|O SߠO�O�O�O�O�OO _0_B_T_f_x_�__ �_�_�_�_�_o�_,o >oPoboto�oo�o�o �o�o�o�o:L ^p��#��� � ���6�H�Z�l� ~�����1�Ə؏��� � ���D�V�h�z��� ��-�ԟ���
�� .���R�d�v������� ;�Я�����*��� N�`�r����������@�����@������	��+�=��,)�n�!ߒ�y϶� �ϯ������"�	�F� -�j�|�cߠ߇����� ��������B�T�;� x�_���O������ ��,�;�P�b�t��� ������K����� (:��^p��� �G�� $6 H�l~���� U��/ /2/D/� h/z/�/�/�/�/�/c/ �/
??.?@?R?�/v? �?�?�?�?�?_?�?O O*O<ONO`O�?�O�O �O�O�O�OmO__&_ 8_J_\_�O�_�_�_�_ �_�_�_��o"o4oFo Xojoq_�o�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t��� �����Ώ������ (�:�L�^�p������ ��ʟܟ� ����6� H�Z�l�~������Ư د������2�D�V� h�z�����-�¿Կ� ��
�ϫ�@�R�d�v� �Ϛ�)Ͼ��������h�*�`,��`���U�g�y�Qߛ߭߇�,���ߑ� ���&�8��\�C�� ��y���������� ��4�F�-�j�Q���u� �����������_ BTfx����� ���,�P bt���9�� �//(/�L/^/p/ �/�/�/�/G/�/�/ ? ?$?6?�/Z?l?~?�? �?�?C?�?�?�?O O 2ODO�?hOzO�O�O�O �OQO�O�O
__._@_ �Od_v_�_�_�_�_�_ __�_oo*o<oNo�_ ro�o�o�o�o�o[o�o &8J\3� ������o�� "�4�F�X�j������ ��ď֏�w���0� B�T�f����������� ҟ������,�>�P� b�t��������ί� 򯁯�(�:�L�^�p� �������ʿܿ� � ��$�6�H�Z�l�~�� �ϴ���������ߝ� 2�D�V�h�zߌ�߰� ��������
��.�@�@R�d�v���qp����qp����������������, 	N�r�Y������� ��������&J \C�g���� ���"4X? |�m����� /�0/B/T/f/x/�/ �/+/�/�/�/�/?? �/>?P?b?t?�?�?'? �?�?�?�?OO(O�? LO^OpO�O�O�O5O�O �O�O __$_�OH_Z_ l_~_�_�_�_C_�_�_ �_o o2o�_Vohozo �o�o�o?o�o�o�o
 .@�odv�� ��M����*� <��`�r��������� ̏�����&�8�J� Q�n���������ȟڟ i����"�4�F�X�� |�������į֯e��� ��0�B�T�f����� ������ҿ�s��� ,�>�P�b��ϘϪ� �������ρ��(�:� L�^�p��ϔߦ߸��� ����}��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� 	�������������
�������5GY1{�g,y�q�� �<#`rY �}�����/ &//J/1/n/U/�/�/ �/�/�/�/�/ݏ"?4? F?X?j?|?���?�?�? �?�?�?O�?0OBOTO fOxO�OO�O�O�O�O �O_�O,_>_P_b_t_ �_�_'_�_�_�_�_o o�_:oLo^opo�o�o #o�o�o�o�o $ �oHZl~��1 ����� ��D� V�h�z�������?�ԏ ���
��.���R�d� v�������;�П��� ��*�<�?`�r��� ��������ޯ��� &�8�J�ٯn������� ��ȿW�����"�4� F�տj�|ώϠϲ��� ��e�����0�B�T� ��xߊߜ߮�����a� ����,�>�P�b��� ���������o�� �(�:�L�^������ ����������}�$ 6HZl����� ���y 2D�VhzQ�|�>Q������ �����,�/./ �/R/9/v/�/o/�/�/ �/�/�/?�/*?<?#? `?G?�?�?}?�?�?�? �?OO�?8OO\OnO M��O�O�O�O�O�O� _"_4_F_X_j_|__ �_�_�_�_�_�_�_o 0oBoTofoxoo�o�o �o�o�o�o�o,> Pbt���� ����(�:�L�^� p�����#���ʏ܏�  ����6�H�Z�l�~� �����Ɵ؟����  ���D�V�h�z����� -�¯ԯ���
���� @�R�d�v��������O п�����*�1�N� `�rτϖϨϺ�I��� ����&�8���\�n� �ߒߤ߶�E������� �"�4�F���j�|�� �����S������� 0�B���f�x������� ����a���,> P��t����� ]�(:L^ �������k  //$/6/H/Z/�~/��/�/�/�/�/�/����+������?'?9=?[?m?G6,YO�?QO�?�?�?�? �?OO@ORO9OvO]O �O�O�O�O�O�O_�O *__N_5_r_�_k_�_ �_�_�_��oo&o8o Jo\ok/�o�o�o�o�o �o�o{o"4FX j�o������ w��0�B�T�f�x� �������ҏ����� �,�>�P�b�t���� ����Ο������(� :�L�^�p�������� ʯܯ� ���$�6�H� Z�l�~������ƿؿ ���ϝ�2�D�V�h� zό�ϰ��������� 
���_@�R�d�v߈� �ߡϾ��������� *��N�`�r���� 7���������&��� J�\�n���������E� ������"4��X j|���A�� �0B�fx ����O��/ /,/>/�b/t/�/�/ �/�/�/]/�/??(? :?L?�/p?�?�?�?�? �?Y?�? OO$O6OHO�ZO�$UI_IN�USER  ����{A��  [O_O_�MENHIST �1L{E � ( �@���'/SOFTP�ART/GENL�INK?curr�ent=menu�page,98,�1�O__0_B_ �y)�O�Eedit�B�MAIN�@RRA�_ESTEIRA �O�_�_�_�37X_j^PEGA_BA�_�o)o;o�>�O�O71 `o�o�o�o�o^opo,23o,>P��1(�o�N148,2T�����_�_�,COLOCeTORNO	2�D�V�as�D55!�����<ˏݏ  ���0�A ����"�4�F�X�j� ��������şן� x���1�C�U�g��� ��������ӯ����� �-�?�Q�c�u���� ����Ͽ�󿂿�)� ;�M�_�qσ�ϧϹ� ��������%�7�I� [�m�ߑߔϵ����� ������3�E�W�i� {������������ ����A�S�e�w��� ��*��������� ��=Oas��� 8���'� 0]o����� ���/#/5/�Y/ k/}/�/�/�/B/�/�/ �/??1?C?�/g?y? �?�?�?�?P?�?�?	O O-O?O�?POuO�O�O �O�O�O^O�O__)_ ;_M_8�O�_�_�_�_ �_�_�Ooo%o7oIo [o�_o�o�o�o�o�o �ozo!3EWi �o������v ��/�A�S�e�w�� ������я�������+�=�O�a�s�^[�$�UI_PANED�ATA 1N������ � 	�}  f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10Ԑ�Őice=TP&�_lines=3�Ԑcolumns�=4Ԑfonܐ4�&_page=d�oubŐ1��\V)�  rim#�L�  ��c�u��������� $�ϯ�گ���;�M� 4�q�X�������˿������%�\V� �� E�  �W<�]���ʟܝ2�����2/�-�ual����_��"�4�F� X�j�ώ�u߲��߫� �������B�)�f��M������3� �E�  Y,� �����*�<�N�`� ����Ϩ��������� i�&8\C� �y�����@�4Xj=�� ��������� / S$/��H/Z/l/~/�/ �/	/�/�/�/�/�/ ? 2??V?=?z?a?�?�? �?�?�?�?
O}�@O ROdOvO�O�O�?�O1/ �O�O__*_<_N_�O r_Y_�_}_�_�_�_�_ �_o&ooJo1ono�o go�oO)O�o�o�o "4�oXj�O�� ����O��0� B�)�f�M��������� �����ݏ��>��o �o���������Ο�� 3��w(�:�L�^�p� ��韦�����ܯï � ���6��Z�A�~��� w�����ؿ�]�o� � 2�D�V�h�z�Ϳ��� ��������
��.ߕ� R�9�v�]ߚ߬ߓ��� �������*��N�`�G����	�������������"�)��G��� 6�s�����������4� ������K2o V���������#�����$U�I_POSTYP�E  �?� 	 /��UQUICKME/N  ds��WRESTORE� 1O�?  ���! /#���m+/T/ f/x/�/�/?/�/�/�/ �/?�/,?>?P?b?t? /�?�?�??�?�?O O(O�?LO^OpO�O�O �OIO�O�O�O __�? _1_C_�O~_�_�_�_ �_i_�_�_o o2o�_ Vohozo�o�oI_So�o �oAo�o.@Rd �����s� ��*�<��oI�[�m� �����̏ޏ����� &�8�J�\�n�������ȟڟ�SCRE��?�uw1sc�u2�U3�4�5�6��7�8��TAT�`� ��MU�SER�����ksT���3��4��5���6��7��8��UN�DO_CFG aPd����UPDX�����No�ne���_INF�O 1Q�<��0%��W���E��� i���������տ� ��:�L�/�pς�eϦ���)�OFFSET' Td@���{� �����	��-�Z�Q� cߐ߇ߙ��ϝ����� �� ��)�V�M�_�q� �۹�����
����t��)�WORK U4�����A�S���ψ�UFRAME�  ���&�RTOL_ABRT���$���ENB����G�RP 1V��?Cz  A� ��+=Oas������U������MSK  �<���mN��%4��%��<)��_EVN������>�2W��
� h��UEV���!td:\e�vent_use3r\-�C7���}�F��SP���spotwel=d�!C6����!�Z/�/ :'�H/~/l/�/�/�/ �/-?�/Q?�/? ?�? D?�?h?z?�?O�?)O �?�?OqO`O�O@ORO �OvO�O_�O�O7_�O�[__Z]W+�2X�����8V_�_�_  �_�_o�_,o>oobo toOo�o�o�o�o�o�o �o:L'p��]����$VA�RS_CONFI��Y�� FP{����|CCRG��\��>�{�t�D.� BH� pk�a��C�� ��}�?�x��C,&Q=��ͩ��A �MR2bN���	}�	���@�%1: SC�130EF2 *(����{�����X� ˂5}�����A@vk�C�F� w�Q�[���|�����������T����\��ϟ �\� B���;�e�@�ǟ`��� ��S�����̯���ۯ �&�}��\�G�Y���pE���ȿ�TCC�Ac
��������p�GF�pgd���-�23456789017�?��ׁ$���4�v�Nm�� ��϶�BW�����i�~}�:�o=LA� څ�6�@�6�ͿZ���$i�7����(��W��� -�]�X�jĈߚߕϳ� ����������%�7� I�r�m�ߨ�ߵ��� �������8�3�E�W� ������}��������� ����/�A�S�e�w��MODE��t ��RSLT e�|k�%"zς�� ;�1��d��`�>�SELEC���c��	IA_WO֗Pf �� }W,		���|���G�P ������RTSYNC�SE� ��$�	#W�INURL ?*ـ�;\/n/�/�/�/�/�uISIONTMOU���A#� ��%�gSۿ��SۥP��� FR:\�#\�DATA\�/ ��� MC6L�OG?   U�D16EX@?\�'� B@ ���2T1���?T1�?�?������ n6  ���GV�2\�� -��5�� �  ��Z�@U0>58TRAINj?��4*B{Rd_Cp��F'#`{2�'$�":��h#� (�kI �Mw��O�O�O�O�O1_ _U_C_]_g_y_�_�_\�_�(STA� i�B�@�?o0oI:$o\bo�%_GE�j#�;�~@ �
�\�|�btgHOMIN�_kSۮ��`�2(,,��CWǖBve�JMPERR 2=l#�
  QoI: ��"�4Fwj| ��������l�&%S_g0RE鰹m�^۴LEXdn��1-ehoVM�PHASE  �e׃BޱOFF� _ENB  ޢ$VP2�$oS�ۯ��x�c C�;�@ �@�;���?Gs33'D*AA���]� ��0ޱ�`r}�XC��܅���\A8-۟E ���� ��#�5��������� ����}��������� �c�X���A�����ϯ �+��߿��M�B� q���xϊϹ���Ϸ� ������7�I�;�m�b� )ߣ�Eߓߡ߳���� �3���W�L�{ߍ��� �����������/� $�6�e�W���c�y��� �����������O� ��?M_q����� ��'9�=7 Is������ /m/%/3/E/s��TD_FILTE:�`s�k �x2�`����/�/�/�/�/ 	??-???Q?�6�/~? �?�?�?�?�?�?�?O� OoiSHIFTM�ENU 1t}<5�%5�~O)�\O�O �O�O�O�O�O�O'_�O _6_o_F_X_�_|_�_��_�_	LIVE�/SNAP�Sv�sfliv���_�{z`ION ҀyU
`bmenu&o�+o�_�o�oV"<E�uZz��4IMO�v����zq�WAITD�INEND  0�ec��b�fOKو'OUT�hSDywTIMdu��o|G�}#�{C�zbx�z�xRELE���ڋxTM�{�d��c_ACT`و���x_DATA �wz���%  OL�OCA_BARRA_TORNO�o<6Ex�RDIS
`E���$XVR�a�x�n�$ZABC_GRP 1yz���� ,�2�̏.MZD��CSC%H�`z���aP@�h�@�IP�b{�'���şן�[�M�PCF_G 1|
'���0�r�8���� �}'��p�s�� 	(���  <�l0  ��~?S��?���?�  5���^��^���e�������¶���C�y�C�K���1w�?��>����	>��>�-�׿�8�������k�rꫠ��������F���ȹ�T�Ǡ�ˠ�Ϡ�Ӡ��ׯ�먗��  ���o���w����� ˩�3������B� �˴2�۰�߰��ù����	��1�?� i˟���ïբ0ۯ���	��`~����_C_YLIND~!�� Р ,(  *.�?ݧ+�h�Oߌ�s� ������ ��(�	�x�-��&�c� �߇�������j�P� ���)��~�_�q���� �2�'��� � &����������&h��I��cA����SPHERE 2�������� ��A�T/A��e ������ /N`=/�a/H/Z/��/��/�/�/�ZZ� ��f