��  	^��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ��!PCOUPLE�,   $�!PPV1CES C G�1�!F0 A> �1	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q�RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Nb_OPT�2 �� ELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1� UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t���MO� �sE 	� [M�s��2�wREV�BILF��1XI� %�R 7 � OD}`j��$NO`M��!b�x�/��"u�� ����4AX��@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC���a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���OR  �BIG�ALLOW� �(KD2�2�@VAaR5�d!�A}#BL[@S � ,KJqM�rH`S�pZ@M_O]�z���CFd X�0GR@��=M�NFLI���;@UIRE�84�"�� SWIT=$/0_uNo`S�"CF_��G� �0WA�RNMxp�d�%`L�I�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�S�� X�r$OR�I�.&ӧRT�`_sSFg�CHGV0I�p�T��PA�I��T��0��>� � �#@a����HDR�B��2B�BJ; �C��3�U4�5�6�7�58�9>� ���x@ޮ2 @� TR�Q��$%f��ր��Ɩ�_U����4@COc <� �����Ȩ3�2��LLEC�M�-�MULTI`V4�"$��A
2FS�GILDD�
1g�Oz@�T_1b  4� STY2�b4�=@�)24�� DԼ� |9$��.p���6�I`�* \�TOt��E��EXT����ї��B�ў22X�0D��@��01b.'�B  �G�Q� �"Q�/%�a��@X�%�?s��E�U� S���;A�Ɨ�M�� �� CՋO�! �L�0a�� X׻pAβ$JOBB�����f���IGO�" d Ӏ�����X�-'x���4G�ҧD2�_M��b�# tӀF� �CNG�AiBA� ϑ�� !���/1��À�0����R0P/p����$
�|��BqF]��
2J]�_RN��C�`J`�e�J?�D/5C�	�ӧ��@{ :��Rd%�������ȯ�qGӨg@NHwANC��$LG5���a2qӐ��ـ��A�p��z�aR��1��0Ex�>$FDB�E3RA�cEAZt@��ELT���в`FCT���F࠳`��SM� �I�lA� f��f��&��5�5Є���S[�g���M`�0��`���#HK��CAEs@͐��W���N���1CpXYZWH�`�����&	��d����&�2�!SWAq��"��'p�STD_�C�t�!W��USTJڒU�()�0U0�!%E�1�!�_Up�qn�) \�1UM)1ORzs>2p;���`YO< RSY�G�  �qd5Up��H`G���{@�c�%0PXWOR�K�*0�$SKcP_�pAq1�DB��TR�p + ��C �`����`m�U DJ�dp�_C"�;b�3 �7PL:c�a�tő"��D�AGQ92����Q�PV.��DBd��,�2&1PR'��
_�DJa9��g- /�P�$r�$Z��L{I.L�Oz�����/�O��CPC�0�O���r~�EM�c� 1�O��C\@RE4��B2�H $C)b-$L>S.${Cނ��O[INE�]1_D!V`ROyp�������q�S=�z0�VPA4���Rp`RN�R��MMR(�U��I�C�RmPEWM0�SIGNZ�A����U�a/$P-�g0$P�s�1`B�`-ds�1`DIp� �-�hTTQ/b�GO_AW���0ؑ�H!$0CSd�.�C%YO�3���P1}��a�vIG2�j2vN��}��K�c�cO�4� P $��RB,���PI�gPKwq#BY��p(wT=A�d�HNDG�A5 �H4��!wE��%�$DSBLI��us��fm0��y@�aL۱a6Url0]��xFB�|�FExQ>��r�d�c5��7D�i�Z!���MCS��pl4&��ra"H�W�K������L���O��aSL�AVQ8��IN�P^�(v]����a��9/P + �S� � �~�0 �0��FI2����烤-1�r-1Wr��NTV��rVݑ��SKI�TE`5g�@��Z!�J�#@#_�@j�SAqFT�a|�_SV��EXCLU��T0JpD\0Lr�Y�t<��Y�HI_V b"PPLY@6�ёS����ӓ_MLs�T0?$VRFY_�3ђ�M��IOC�[�C!_��2��Op֕�LS� |rLD4$A$W��c�о0P�5,�l�`)�AU��NFzv����e���`s�:1CH�D��up������AF�I�CPr�T$A8����q :P�0qT��� z� �ds_N��c� ;����T��� ��E�����SGN��<A 
$ �P�QdQ��o�9���0#��2s��2��ANNUN�@�����e IT0`5�˹ȱ�Xк�"2EFi0I�B=v�$F��4 OT�P��LDj�NB2Ahb�IA�M�pNI�B!>��Z��\�A��x��DAYC3LOADЀ�ADS�MC5IA_�EFF_AXI�r%?P7AU#O���C��0_RTRQ��@� DWp/P��Q�"B��E|`�ø���?��`�� ������MPE�� A\�6���06�Jc��DU�P��]��2CAB��B�fPNSH���ID��CWR �3�\�Vw�V_2������DI����$C� 1$-V�PSEs�TW�p��M���$@dE�_��J�VE�� SW��a ����d����@ ��OH��fO�PP�K�IR1B�0��Lӥ��R�! 氃�}#}���}�v�s��B�����`��R7QDWl�MS} ���AXR��J�LIFAE�0��SA�N� (�ȱ�C�wǳ-CH raN*�z�R��ȱOV 4�H�Ew�SUPPO$�0{q��0_��y�BW�_���ma��Z��W��H!���ȱfrq"cXZerA��Y2EC_PT�0�P��N�T��ȱJ� d�_�����YA�$D =`�`CACHR����SIZN�z�b�� SUFFI������0N�AD��MC6�IA�Mv vE 8�԰KEYIMAG�STMRQ\�Q�����2W�OCVIE$)�01F�"�L!�n�^ރ?� 	��D�jvG��@�STM�!i$@q2@q���q��qEMAIL�q��P��n�ءFAU�L�BH�"�S�3AXby`U� �P�@DT-P~�!I< $���S2Г�IT}sBUF�ށ��d00%��B$tC݄ԡ8�3�SAVS%"���:�3�n'��̶P Z$�0P*�tp_ 9%�r��)OT�R��ңP`�:@�*��'AXC3�	��X z��#_G:�
n�YN_t�J <WpDuA@�uUs�M^�n�Tr��F�P$�P��DIB��E�0-P.��1K�ǐG)!$�&m�jQ`1�m�p�Fyp L (PSVw`�dADM�6�y[1�2�Q3Q�M�:P�1��#C	_�P�PK�T @���4�w�R��5��1DS�P�2PCAKIM@`#8C^Aߥ�1��UG0��U ��IP"��3]�Y 7DTH9 �s+B2��T�Q8CHSk3CGBSC/�H PV����J�@�#�DD`��NV���GS�D9 5F F�� 0dC[0�!�QSqC��u�3MER̔>yAFBCMP̓�0�ETa� N�FU��DU�v��PڒCD.I�@� ��PQR-���c�O���`��Rr��T��P,��RC"H��U0�2U�S|� �PH *�QL����a�!cV�b� M�Yd��WfH�Wf��WfP��Wf�Wf7Ti8Ti�9Tj�Vh`j1mj1�zj1�j1�j1�j1��j1�j1�j2�j2T`kmj2zj2�j2�jU2�j2�j2�j2�j�3�j3`j3mkzj3��j3�j3�j3�j3ʻj3�j4�b�EX	T��c�Q22�70K��70QeB0���U����FDR��RT�V}��"����B.�REM�Fla�ҧOVMC�A�T7ROV�DT^ /�MX>�IN�`�.�N��INDM�
y�l0 050G1��8�_�(��D��8�RIVx��L���GEARAKIO�K��N[0�호��*��� Z�_MCM ���F��UR�RS ,<�Q+!? _�s@s?K��?K��EV�S�mE!oPՂT� ��P�!��R�I�p�#ETUP?2_ U ��##TD�@V�$T��c�p����H���BAC,2GV Tj����4)�:�%�cV0�PIFI�`�V0oP@`��PT�+��QFLUI\�W Щ�>�UR ��>!f�"s1�@ �Ӫ�I�$��S;�k?x��J�0CO� ��#VRT��%�x$�SHO�װ�AS�S�@�!N��@��BG_�s�
��zc鱇c�鱔cFORC�_^D�DATA��X�KFU6�1`29�2`1p�E�9 ��Y |��wNAV� ���ʷ����S�L�$�VISI�� bSCF�$SEq�Ӱ]�V��-O��$�PB"�`��gй�$PO��I�k��FMR2>҅Z ߂�P �����0�������P&�������_�a����IT_5��T �M���ɟ۝DGCLF�a�DGDY��LD�c���50���(�́M��`^[%R� �T�FS� ]\ �P��.�3 0$E#X_.�E�.�1� 4P�k�/�3g�5g��G�Q��] �c��RS�W<%O��DEBU1G���GR �UVSBKUaPO1n)p -�PO6Р�����P����MҰL�OO�#�SMb�E�b"��k�L�_E �^ ؤTER�M7�_@��PORI�y1<�`Y�_�SM�_�0��<�aY�J�A�~�b@���UP3c�� -j���^(��N���_��G����/ELTO�d2PFIG�e16����P|e���`$UFR��$�P��) �Um�3OT6PTA�@���HNSTz0PATx�A� ^PTHJ�QҫPE_�3��AR�T{ ����{!�d1R�EL�
�1SHFTP�Be1d�_��R�P��S}� ��$��� b���ဲ�sC2SHI�� ��UPb u!AYLO�@1&1H�t�ɲpdY��U�@ERV_` /}����Dz0��q0'��
�'�RCs��U�ASYMY1�Ue1WJ���E����}��QU�z0&1��Є~�PqCL!QOeRz0M�À�GR&���d4����c # 1敠HO#��e ԰J+����POC��|���$OP��AAEcճ�����0���� R5S�1OU,�Cdem�Rb�%��(��4e$PWRf��IM�%`R_�#`���~�we1UD��ty$y4f��$H�5�!q0ADDR��H�)�Gf�11x1��R�R��2ag H��S \P���s�5
��5zc�5ƇcSEVѧ��PHS<�P��h $6�� �_D����ɲ�2PR�M_i�x�HTT�P_�PH2ai (��POBJ��x2�$��LEUz 4A3`�j � ��yQAKB_z�T�BSp ��CW�KRL'9HITCOU�D갟 �� � �B����ų� )�� �SS~�RdJQUE?RY_FLA��yQ�B_WEBSOC����HW�a��2ak��0 INCPU{��OEV�A_d\R�4�]Q�4]Q�b��IO�LN�l 8��R��{�$SL��$INPUT_,��$� �XP�� �G�PSLA�� m�P�_�U�T��U�x!IO@F_AuS�n�$L�ZG����92`�0�S��S1HY��ca�<c��Q_UOP�o `(`�a��]� Sd]�Zf�a� P=3� ��g�aZf�b�f�1IP�_ME��M�p X�(`IP0{�r_N#ET{�P���"��8"vŁ��DSP�,@��ްBG{�B���M��M�q lM�TiAGa@A#�TI�e`
%= 6Ѝu� PS�vBU6�IDZмB#���u� �ux�[r�rV �r�Rmz�t�t�PN� �6���IRCA|�� s �xIm�PCY�0EAKc�B���G�]�=3_���R�~ ��s!DAY_<�p�xNTVA\��pࣇ�R��s��SCA�A��CLڑ�qɱ��r��M�t�����N_� C-� ��r��N�u�R+��#S��a�UB�p�q@��+� 2t �P\q�M��v��UB�pLABpV��6Ю�UNI/�9��h�ITY�c\q$�5bR ��w�Rd��R_URLk��$AL�EN������t~�ST��T_U�����JDPM�x�`!$;����DPR�e\�"t�A���Qf�J��r�#FLP�4��
�����
�UJR��y �x@FX���"���D��$J7@O^�$J8ܩ7��H�����7��ؠ8��ۡAPHI��Q��+�DB�J7J8�ɲD�L_KEِ � �KPLM�
� z <�X�R`RPȳWATCH_VA��L�QFOFIELpu3yy�L`���{ i�LVU�7���CT
�̶u� �LG��|�� !4�LG_SIZ�D�����`�FD�I�"��� 
�9��	��#Ä�� ��`��9���9��ƪ8������_CM:��W���D�F�����	�r�$(����"��"�`"�9�.�I�!�8��"�9�"�	�RyS��s   (��SLNС��}�`�@ ��W��RO����C��rp L�Ӯ�DAU�ՃEA#@P�$����GqH�"�+`BOO�1?~� CBb70�ITS� >fREbp5�SCR
ЪCCa�DI=cS# �0RGI,�$Di��V6c�$H���D+aSfC*bWq�+a��6cJGM��MgNCHS+aFNV�b��K��$���UF�����FWD��HL.5�STP��V��ԐX��%���RSm�H& �3fCK��6cT ����UA���:ӳ��ְKc�G�� PO 	P�`�K�����Nq ��EX2gTUI��I i�9�>�i��~�� ��ّ� ��:�	؀R��� Q�NO�ANA+b�!��AI�D��DCS���3�3*O
OSy�4r!S-��IGN"����4����b�DEmV��LL�G��s�`���qT$��$��MR8���K�Ag1���	��PXS\q� OS1�2�3�   ��`G� �xK���U 4�T�uAU$ 3���Vh&ST�`R��Yp�� �  �$E�&C�+Р@�&�&\�9�a� L?PQo��`fh'v�#�@97EN#@�;4
�O�_ � �@��)@ՃR�J3��MC��� ����CLDP�`N�TRQLIґP�~9l4�FLSq�2A�3�D���70PLD�5�4�5�ORGV���2��RESERV`T�4lS��4wR ]3��� �� 	�5��{4�5S�V��~0��	�1YD>aFRCLMCoD�?�O�I�PaA �MDB�Ga���m�$DEBUGMASTc(��~���U��T� �u�E��q �MF�RQ��� � ���HRS_RU��Q1U�Ac���FgREQ�'�$� �OVER�p4�pt6&��P�EFI�p%�!V��A5�R,Dǈ \F�?Q��$9U< S�?6@��SPS�q�	JSC�АpC|r�S�CU��A�?( 	��MIS�C��� d��<!R5Qo�	@pTB|��pc 3f�@hAXs2�[�Cg\lEXCESH�!bM�`����p�'bs4@ cS}C=  � HP�7d_��1hf��kZolh
�@K����Rݢ|��E{B_ްFLIC�$}B?�QUIRE��MO&|O6{�V[1L:0M��� D0-��sp�soB$AND�џ�����Ҡ����s�D�ü�INAUTb��RSMѠ�xY�NRB����q�A�qPwSTL��� 4�7LOC?&RIԐ?%;EX4�ANG��RkL���AU�#`1����L�MF�@� qVe)2��5�����FgSUP(6	PFXi��IGG1� � �6@3��V�3��4 �R�"牌 ��� �`�`&~���QTI����`��MY��B� Mtg�MDd�Ȓ)r�
}��Az�HH��}�GDIA�~�l�W��P}���}�D��)�aqO��W@��� �`�CU"�V��Q@�Q�ʧPO��_�@��� ����G#q��@�R��D�.�P.�x��5�P�-�KE���-$qBYP!�� ND2�B���~�2_TX4XGTRA
���B�spLO�з���b��/b���Җ���أ�rRR2e��� -С��A^A ?d$CALI9`���G��2�RIN�� �<$R*�SWq0�DZ��CABCx��D_J��-q�q�_�J3��
�1SPHް& �P���3��(��� �յJ�C�4 BVAO�IM�@�RCSKP�:�����J���RQ�E�+�8E�;�=�_AZ]B��w�EL�ಈAOC�MPK� a�Q��RT�A��ҥ1����=`�1��ȩ ��Z��ScMG��U��DJG<0�SCL|`8�SPH�_9�Pe�Ӗ���'�RTERY� ��� �_� K1d A0���#�RU�DI��ҷ23U�DF vv�LW|�VEL~1�IN2� ��_BL 
�R����QJ�Ԭ�<�׽�L�IN8�?Q�`����Ջ����� _` ����]Ո]��b��m� D�H|`���a��$aV)��sө$��XUQ0Ro�$���P�R蓶`�H ��$BEL��W5�_oACCE�� ��<�A��IRC_V�p���0NT�Qi#$SPS|`q2L <� ��3����m�� ��u���6���6�3��a_���g�m�PU�P��7_MG/SDD��V�0RFWa0V����������DE��PPA�BN�RO�EE }����~0;���A�`��� $USE_t(��PYPCTR��Y���\A �!YN�`A� T���TM�A ����O��(�INCڔE����@b���AaENCF�L�<��R����>d��IN�q"I��W��NT|�Ӿ�NT23_z�0RLO��0R.gPI�pO�9��0c�@8��0��bC��MOSI���b�m�OS�RPERCH  UeQ;� �K���; �D��Ǖ�>D�l��	A��L4��g�� ��;6&QTRK9�1AYԣ��af! �u%j#F����a�PMOM�@b�b�0��/d����#8���DU
�b�S_BC?KLSH_C��% �@vfP\�S3�!:|k=�CLALM�p�A� <�S5CHK�|H���GLRTY"� o��I��1U�_��k'_UM�C�6C�C��Ѿ33PLMT��_AL�0���4���7E�= �0�;�0���5�跰�C� ">D�PC��HpTp���5CMC��\���CN_7�N��L�F�SF���V>�G��5�rA��EvHCAT�>SH��7��� ��1�!�ѥ�ѩ��f��PA�4�_P�5�#_��m&��}#�T�5JGx��`�S���OG�GA�TORQU0 ��i�)��r�B����R_W�%f$��@��d|�e��eIkI(kI��F^�a�Xgh����VC��0�a�e�b1�n��o^��f�JRK�l�b�f�D�B
�M&��M�p_sDL|�"GRVd`t|�t���aH_ף8�c9�@zCOSM{��MxLN�`p{�ewt|� ry��ryDa�z�|ba�e1Zkp��aMYyq�x�Yrw�a{�THET=0N�NK23��7�lv�zpCB<�CBv�C,�AS=�a�Ddo�|�o�<�SB|㍂G�'GTS�C��iQ���XS��Ê�s$DU}0'��������eQ�_RC*QNE�%�K�4��[�Z�+��A/�X�a�?uJxJqLCPHMu6�6�S�e ���u���u6��vӓ���vX�Vz�Vo�l���UV��V��V��VʛUV؛V�V��Hz�@������Q����H��UHʛH؛H�H���Ok�Oz�O%���O���O��O��OʛO*؛O�O�vF6�\�𸹜u��m�SPBA?LANCE_�q��LE��H_/�SP��эvv«vPFULC�;�#�;«u���1���UTO_<x0�5T1T2|ɼ�2N_1�������!�=����!T' O�o���`INSEG��ZREV��Z�gDIFP%"�1��6m�1�OB��C1�s�'2�Pj1�dL�CHWAR��q�A�B_Q�%$MEC�He��psyю6AX�s!P!D��Q�]�q��� 
���Q���RO�B�CR��ՇB ��C��_{RT� � x $�WEIGHp A �$k��PIp6I9F(��LAGa@BqSa��aBILG�cOD� ]%�ST��"%�P��C0&��� P���О�
� ��b�{Q  2�h*�D�EBU6�L.�v���MMY9����N8IS��A $D.��$���P� ���DO_��A�џ <�����1bN�IB`�X�N�3�_?�b  }�OP0 �/� %�0T� ���1T������TICYK7�K�T1 �%��� ��N�k�'�R�0b[ң�[ү��P�ROMPpEM� $IR�P`�08��
 )MAI�`�4r_A�
�t|!t RpCOD��sFUh 3�ID_��E�����G_SU;FFD` ;�W
��DO������Z��GRA�[҃�� �[Қ[Ҧ�Q������H1�_FIv��9�ORD`�3 ���36%B�|` �$ZDTL��}�
��4 *	�L_NA<��S>��DEF_IcS ��o��g��q��������IS��@�.������m�A��4�A8Bq�Do��"$ʕ�D�PO��LOCKEIQ}��������} UM�S� �������#� ~���o��&�� f�|Q�S����')5V�P/��f���4���Wd(c5Z#����TEN1��� ;�LOM�B_}2�70%�VI]S[pITY%�A�Q}Oa�A_FRIlÌ�30�SI��1 �R����7���73��%�WB�8W�;p�6�`_4I�EAS-��Q�4P.P* 	�64�95�9�6.�ORMULA�_IIQ�GC�� h ��7��C?OEFF_Ou���H�Du�G!Q-�S6����CA=�����}�G�R� � � �$Z ��(�Xe�TMM'ETZ%{�b#_\1�ER��TC$B� ��  e�LL�" S�M�_SV$�X$Ć6� �аD� � �7RSETU�MEA��b �`&�}��>�Х � �P�� ��@a��a2!D)fX��2!N!/$�RA�Yc��+ ��* ek�2� R�EC#a��MS�K_�+S� P~�1_USER������dJ��t�`��VE�L\b�`J��b�e[�I�,���MTV�CF}G�a�  ��z�O��NORE���;�r�K�r� �4 c|�3��XYZ���������3po_ERR�ѩ ��PT�5 Szp��`��`��BUFIN�DXOa�0��MORn+T� H�CUzq ;���q+�c���O$���v��Nb�1���G-R� ?� $SI�@@5 ���`VO(�#����OBJE.�)�ADcJU��+�:�AYWP4��2�Dh�OU� Su��pa�=�qT������`��
�DIR�����
������DY�N&B��߅Tp�S�R��1f�`�R��OPW�OR9� �,>��SYSBUH�Pa�SOP!��r�Q,�U�+�
�PZ �bR�PA`�`#aT�}�PaOP� UR�F�/ђ��Ⴠ/IMAG�q���fq�IM�q��IN4@�z���RGOVRDԁC��`��P�����Р��0#����LX B�wp��aPMC_E(4�q��NH�M$���b��1��`ԑSL.��`� ��OVSuL��SX2DEX!D�i�2�����A_Ԑ ��� Ր��� ����������C��U��ϡ��^Ր_ZERqH��S�a� @@p좜�MOM RI+���
�� �2�%�q�E�Lʭa��rT~�u�ATsUS`��C_T���rm�BIPw�`�"d#p��L�4�`� D� ��l�j�ܰ��k�����a��XEq�*eŲٲĤ���	��p�UPXd��PX�𗶀����36�����PG�u��$SUB�_����!_�3�JMP�WAIT���w�L�OWMs|�)�E�CV!F����z�R��p��CCҠRց����IGNR_PL3�/DBTBu�P���#BW1 ��&pUH���IGj���I��TNLN���R�S"�0yN��c�PEED�>r�HADOWu���&p3�Eq�kԀ�I�nwSPD�a� L��A��o��M���UN�#�:˗��R�ڣL�Y)��i��P�P�H_PK5u�rRETRIE3�*r���$Q����FI8r�� �X���� 2}�pDBGLV��?LOGSIZ,�!KKT��U�SP�DV�n�_TX�EM�@!C�ad�v�_�Rp�L2>IvCHECK
�Oa��P�`�Ѷ�p�鿂LE"�RPPA�A T��a�ms��P4Ҏѷ�BARC�8Ӱ��E�O� Nr�@ATT�ҖaC�v�0)b!.��UX��r��LJ t� $q~M1SWITCHr�ZQW6�AS3����q�LLB�ѹ�_ $BA�`D(#PaBAM�ă��3����J5jp q��6|����_KNOW��4ԀU[cAD��P��D�`%	PAYL#OA#a� C_�qLT$�LZIL�!AaާLCL_�p !�P����a���F�	C�P�
"b��@I�R�P��r��BU@�qJc�
_�J��a�qAND��rsb(����@AP�L��AL_ �@~���p����0C\buDHE[b�J3=�Q� T�@PDC�K��PaCO�P_�ALPHa�BE0�q�Aas �
R�>� � �L�BWD_1I
2sD�PAṞ$(%5& #��TIA4O)5O)6\bMOM�p[#{#h#h{#u#pB��AD[#p�&h#�&u#PUB�R�$�%h#�%u"��r���d�� L$PI֤2� #�aN9ɡTh	9I*;I8;IF3�, mq�w6-�w68������s���O�HIG��Oӏň��6�ԏ� �����6�3�8���9����SAMP԰�v2D��73C����.  �PaA�pq��rpD-�zF �� �I  �r���X �xEM��H �zCIN �LMC�H�K�D���J�
X�D
[*[GAMM�ESs�_t$GE�T�2�pQ�D��b
�$TIBR�0�I.jw$HIX`_đ�p$�r�VE�p�XA�^�P�VLW�]�V�\�Yf��V��6&�SC��C�HK���`�I_@���tL�L�E�tg�#�t�&siQ ��$� 1�� �I1�RCH_D����RN��V��bLE���2� x��`}�3�MSWFL���MQSCR"�75��L�pD3W�Tv�G�p�[ �Ihy��wt	�#SV�ѾPـ��;wίqGROU��S_�SA�����u�NO�C����p}T� TfL8:�*�r0z5,g� #DO��AzR�� qEjz�E�8&��6���80ˇǅ��� ��q�}M�%� � yc#YL3��GGPL� �W����%�	��d�)����;p��ñM_	W�pk�q�� i��b��M����� ��P��A:�q�9�-�� M�q� 2� �!����$Wݐ`�ANGL F�vݐ�ے�ے�ےu���PN��S��q�MX��O�LZpa�� ���$� �,aOM�c��!�3��E�W�R ��b���L:�_x�� |��� �p{)'�h#'�u#�pT* T�?�n*��wU��
��r���w �P��PMON_QU7@� � 8��QCsOU�aY�QTH�sHO�ҰHYS4�3ES��ҰUE���r���Ov��  ��P����U�qRUN_T�OI����2�p� �P? ŭůqIND9Ep�� GRA��h��*�2q�NE_NO�f��IT�`h���INFO�q���Nˏ��(�������� =(�`SLEQ�6��0�5��R�ِOSM`���� 4��ENA�B	��PTION�(�k�2����GC]F�� @��J��,L#���PRK�����,��"EDITN�q� �!�b�K�j�3�QE�PNU��Ξ�AUT�q��CO�PY�ѭ0�܍1�pM�QN����EfPRU�T� ��N=�OU���$G �+��R�GADJ����X_r�I�c`�W�n�W�WU�PU�pW��3G�z�RN8_CYC	����RGNS��͜�@LGORc�NYQ_FREQ�"AW�@�6��B��L~ �*���U�v#�@�5CR1E�PݳS`IF81Z��NA;A%&�_G>�cSTATU��c��MAIL9BI<qʹLASTq�޺�ELEM��� ��5�FEASI �˂fB^pQp��1�q��ҭ@�PIs��d��`�1ձ��sAB�sE_��0V��
�*	�R�!U�0�0�p�SRMS_TR L�`nY��0�R���R �����#���	�� 2� �CF��D�� ����@M��7�d'DOUH��dN/Ӽ��PR�������GR�IDm��BARSF�7TYӵ��@O� ���� �_B�!ȃ�i)O_���� � q���PORpHÒ6�SRVF�Y)��DI�pT @���0��0�4�TKp�6�7�8�Ҵ�FZR���
�$VALU9�u��|G!���� ! Ո��\�|H�x�AN�sp"X�R������TOTAL8C<��#�PW��I1�$REGGEN�*�"�X_`0��噱�&��TRE�2�!_S�pE7� �AVU�p�f2.�Ex��5ױ��¸Ъ#V_�HRDA��e0�0S�_Y�qY���SFpA�R��2� #�IG_SE��O0����_��4C_]$C�MP��BDE ��0BIUaZC�3�Q�CG!ENHANC���� p��8X�S�1INT��!�F�}�MASK\T�P OVRݳP�� 5ԠG�aF�E#4����B��;]�P�SLG�0���C�@�r��Qr��� � SX���!AUPqƶ��PTEQ�P ���� �QEeJ�F�r	�IL_M��Pso0��TQ���Cr�Y wL�5V�[C�]P_�P�p��SM�YV1�ZV1��[2	k2�[3	k3
�[4	k4�Z�qk0kr`�q.ІfZ�lrIN�iVIBȐ�T�`���dU2�h2�h3�h3�h4�h4�h���RQ�r����T $MgC_F۰�p���L�q�qaE� M�pIaC>r
 ���!B�o�KEEP_HNADD7q!yt# �y	C��F��ti8r+P�sO��xt�6qn0�s\fG�sREM�r�t��!��u�q�xUB�e��tHPWD  �ysSBM�A�COLLAB���  P4�!,���IT��P����NO��FCAL� �u}�� ,��F�L�I$SYNT0p��M��C�2�� �UP_DLY���
�DELAɀ�!U�Y��AD���AQ�SKIPߕ� �4��O+�NT�aM��P_�F��N�E� � )�k17�.�7��6�  6� 6�& 6�3 6��@ 6�9��J2RT�������XD T�� ؑ����ؑD�urؑm��uq��RDC�!��+ ���RL�R���P��aR�"�ղ!��R�GEY���)�FL�G����9�W��SsPC�ç�UM_ؐ�wS2TH2N���ː 1� ��ːi�� �� D;�[Hq�' 2_PC���SIQn���_L10_C�pܼ��A �O�$ 젘���*���R�Q+�)���hѪa��)� b�]��"�2't!��t@*Ǡ�9�D�G��VL1�1�����;10�p_DS�Qq�~�5��11��� �ljp�q<R�p�]�AT�p,���'�R�V�������PҞbHO�MEH� �2������"�4�F�X���3���{ύϟ�P��������4������
��.�@�R� 
�5���u߇ߙ߫�L���� 	��6�������(�:�L�^�7���o���������8���������"�4�F� ��FP�S=�v��  @��0m���pE�� T͠���&��IOtQ	I���2Oy�_OP*B�"l��j�POWE�a�# �����¾$� 푅y$DSB!PGNA���#Ā�C��r!��S232N� ��n��p�HPICEUS�#S�PE��i!PARI9T�1�!OPBe�h"oFLOW�0TR��4�"�qU�3CU� J��j!UXT�Ai!t@EORFAC��pU� ���SCH�� tjp3p_� @w�3$�0�0OM�02S�AR�7�/@9qUPD�Pp
�{�PT��EE�X���nPEFA�Sp B�1M#� Hсh@�" �SZ" �a����qK!  2�� �S�w��	� �$��م���c%?#� _�0J&D;SPV&JOGt0���n�N͐ۅ����6K�_MIR�r!�$�@MT�S�#A�P�S�@��� D��S��0� .���@�%BR�KHi���AXI��  2�C2A"��A�2?#� BSOC�J&�pNF5D�0Y1�6s�$SV�pDIEG�F�GpD��D�B�#OR�7��N�^@�6F0�7o OV�r%SF�:�0�3�BFx�6/�#UFRA�:;TOLCHǂۅV�POV�En!WE�@K�o#�q�2S0�_�0�]� @|�TINsVE[ ��OFSp@C��SWD�13D�1�R1z��%l0TR��<��u�E_FD��!OMB_Ck��BB�B�P>����B�AS�y0�V�q�R�:�ك�2G�G�(AM�#�@jUZB5__M�@/s��g@T$	�)P���T�$HBK��&�QI�O���U:�QPPA�Z�Q�Y�T�U@U:~gBDVC_DB3� ���P���PK�/	e�`hZS	e3f`@Y���?� �1U��d CAB����@L�h�@X��O(PUX�&?SUBCPU�| S1�C��T�C��i��CTv�$HW_C���C��P�fS�q���p��$Ud��#4ppATTRqI|�*r| CYCԢ�{aCAVb�#FLT?R_2_FI��	�\c��P�+CHK�+�_SCT�#F_�wF_ |�r2zFS8��BrCHA1��wp�q�B$�rRSD��`�31��: _TX0v�B`�CEM����EM3T�rC���r��_�DIAG�R�AILAC�S�bM�( LO60��\6��'$PSb"�� p`e�,cPR�PS��]��ǂC�Q� 	YCFUuN�>RINE������r��0�S_����lP��zT�d�zTCBL��&�B�aA;�7q>�7�DA!00�|�B�;�LD�t0��Q��W!�����T�I��ĕ&A�$C�E_RIAu��AF�`P��R@���T2��C�.b�AOyI�p�FDF_L��X�2��LM�CFr��HRDYO�!z@RG��H��!����C�MULSE3��c�g]3�$J�:J�2��7�;FAN_AL�M��¢WRNʥHGARD��n�PqB�2¡�q�%_.@��&AU�@R�t0TO_SBR:/�c �7�p�S��O�MPINFe@,qb���m�7REG��NV�z�j6DU N�DFLu�$M���ptĦd,`h�ѨصCM�P3NFAqxcON�@qж�@|@v����$Ψ�$Y$�&"!+ �� ���#EG��?#t0O�ARQ \52��[�h���%AXEY'ROBnV*REDV&WR@@21_��83SY0��t0��S��WRI@@b��`ST� W#10
�0Eq��k�e3�B_ B�fA!֤�DFP�OTO}���R@ARYV#XҒ�Fd�� �FI� �#$LI�NK2�GTHw���T_�fAj�6�f2��XYZ���7N��OFFn@w���J��\�BT ݂��0CA� ���FIEp��?�l4݂n$_J ���2�ӝQ�0�:ہ8f2� (�Nၢ��CLZ�%DU�ri�9��TURŠX˓��f�b]�X��tPn�FL���@uc\������30�f2|A 1�L�K{ M�$\53�a���e8���g�ORQ:�c! ���a��� O������P���ca!����OV	E��$�M]��#��� )���/���s��wa��p��AN�az����� +���  .b��������L)�L��c!ER�!�	��E@@P���A8h��	�5�0d׃��f��AXCC� ��F`�ay��e��	�� �	e0�
���
���
�� �
��
���
1�� C��	C��	C�C� C�,C�<C�LC�\�C�l�}DEBU�c$���i�-!�B���AB���Q�1��VvP�b 
H"c+� p%�a|'r�|'e1|'�� |'��|'��|'�|'���������y���LAB��n��`�SGROhopn��_PB_C� qԢ3�4�%6Y1o�8U5"�a6AND+�`@`a�Ղ"��7 _Q���в8E��8bp��NqTՠ7C�0VELI���1���6�SERsVE�0>�� $����A�q!"@PO�uB@R�)A��$���ASS  ����PAN�N� }E@VERSIT��NG[@0��aAImp�pNO`@AA{VMՠK 2 �E� ?0  �5WA�Or�H�O�M �LA	P])_N��@�_T_;VYU\x]�_Q`�_�_�_�T�@BS���:� 1nI� <�_o0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2��R@MAXo��5���c  dG�I�NP�b�F�PRE_EXEs�����E��kL��A�@IOCNYV��t� �^�PǦp��s��W�SIO_̠� 1�KP@ ��?Q*��\'��@?� 5���J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_��_�_�_oo0mG�L�ARMRECOV� ��Y����L�MDG ���8�LM_IF �c�5��o�o !z�oDVhz�}?, 
 ���/r;�����!�$ �E�,�i�(�������ÏՏ@�NGTOL�  �� 	 �A   ��G�P�PINFO �k �fP�b�t���Y�  �r����wb ��ߟɟ����9�#� ]�G�m���ġ�ݏ�� ѯ�����+�=�O��a�s������jPPL�ICATION �?������Hand�lingTool� � 
V9.?30P/04���
88340����F0 ��202������7DF�3�����None���FRA�� �6=ͯ�_ACoTIVE=b  ȳ��  ��UTOMOD���u����CHGAPONL��� �OUPL�ED 1�i� �B�F�X�j߼�CU�REQ 1	�k � Tt�t�t�	�����̰��xb�tҤ׵���H��E���HTTHKY��yb�߹��� ��C�U�g������ ��������	��-�?� Q�c������������� ����);M_ �������� %7I[� �������/ !/3/E/W/�/{/�/�/ �/�/�/�/�/??/? A?S?�?w?�?�?�?�? �?�?�?OO+O=OOO �OsO�O�O�O�O�O�O �O__'_9_K_�_o_ �_�_�_�_�_�_�_�_ o#o5oGo�oko}o�o �o�o�o�o�o�o 1C�gy�����܆�TO������DO_CLEAN�|��I�NM  �� tߗ�����͏�ߏz�DSPDRY�RP���HI��s�@ ��K�]�o����������ɟ۟����#���MAX��0��q��!�A��X0�@�=�@���PL�UGG0�1�=���P�RC�Bq�u��:�,���O����SEGF	�K���� q���K�]�o�����˯��LAP(�;���� ����/�A�S�e�w���ϛϭϿ��TOT�ALc����USE+NU(�5� ����҆�RGDISPWMMC�h�C�&S�@@�5�O&�H���1�_STRI�NG 1
�
��M��S���
��_ITEM1��  n�ͼ����� ����(�:�L�^�p� ����������� ���I/O S�IGNAL���Tryout M�ode��Inp�R�Simulat{ed��Outd�OVERR%�� = 100��In cyclX����Prog A�born��N�S�tatus��	H�eartbeat���MH Fauyl����Aler�� %�%7I[m8��� ,��� ,��߸*<N `r��������//&/8/J/�WOR��ۂ!�\/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�?�?8�?�? NPO���� &@�+OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_!BDEV)N�P=O�_�_ oo'o9oKo]ooo�o �o�o�o�o�o�o�o�#5GPALT �nq�/H���� ����&�8�J�\� n���������ȏڏ\GRIF������ :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~� ���R��� *���ޯ���&�8� J�\�n���������ȿ�ڿ����"Ϥ�PREGr~[�ί4ςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ����(��$ARG_�� D ?	����	�� � 	$(�	+[�]��(�>����SBN_CONGFIG7�	�\�[��u�V�CII_S?AVE  (�~��q���TCELLSETUP 	��%  OME_I�O(�(�%MOV�_H������REP���'���UTOBA�CK��	�x��FRA:\H� �2�H�~�'`���H�{�� ��w�� 24/0�6/05 11:_02:20H�?��H�����'l��� Gn�����H��\�,>P �t������ k//(/:/L/^/� �/�/�/�/�/�/�/Ġׁ  g�_J�_\�ATBCKCTL.TM�-???Q?c?\u?<�INIqp���n��G�MESSA�G���1~��;ODGE_D����n��8�O�P�?D�PAUS�:@ !�	� ,,		�?�	�>O LG2OlOVOxOzO�O�O �O�O�O�O _
_D_._�@_z_��D@TSK  !M{��?G��UPDT�0�7d��P�6XWZD_E�NB�4j��VSTAp�5	��U��XIS\�?UNT 2	�{��}�� 	 �o� M7v ����š0b��NH�V`��oXvo�o�n:v��Ġ-hu��Ġ��o�op�o�o03fMET���2�V�� PUa?�Z -?��>��߿4�R�?W0+?^l�}�7GB�7jt��6&ff3`N�7@Ĝ7AUU�9}SCRDCFG� 1	�]� ���{���@�)�;�M�t�H�Q�� �������ӏ���^� ���?�Q�c�u�����0 �:���J�GR=`�PX�?ؓ0NA���s	J�Ֆ_ED�0�1�y� 
 ��%-0EDT-`Ɵ�V�z�Ġ��eP@�K�I�H�?�=x��B���  ���!2�[�8��=w䙦���Ưدn����3 ������d���K� ����:�ȿ�4��� ���)ά��^�p�����5O߿Ϝ���)΀x���*�<���`��6 ��h��)�D������,��7��W�4� {�)��{�����j���B�8��'� K��*̀��G����6���9����*ͨ`Zl��CR� "���X�r�$6��Zؐ%�NO_D�EL�֒GE_U�NUSE�ԔIG�ALLOW 1��   (�*SYSTEM*�s	$SERV�_GR;� @RE�G�%$�#|� N�UM�*�#�-PM�UC uLAY�Op|PMP�AL�05CYC1�0$.7>!0%>]3ULS�v?�%92A�#�Ls?�4BOXO{RI�%CUR_�0~�-PMCNV6��010M>�0T�4DLI�P�?�)	*PROGRA�$PG_MI%>�OOa@AL/EnOXE�a@B�O�.$FLUI_RESU=70�O�/�O�DMR�.� ��b?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o%�7I[6"LAL_?OUT �+�����WD_ABOR�>0g/�sITR_R_TN  ���~�pNONSTO���t p(CE_R�IA_Id �u�0���FCFG� �0��9�_�PA�@GP 1.C�U�����H��Ϗ��C� ���Z�pC��C �(�V@C8�@�H�V�CX�`�h�Up�xꄤ�����R�d�v�l���?��HE �ONFIP���G�_P�01C�  �1#����� �2��D�V�h���KPAU�S�11͕0�  Bj���͕��ܯ¯� ���6�H�.�l�R�|������ƿؿ����r�M~�pNFO 1͕�S� � �	��O�� =��/H�iB9�����{��HџbB/Hl�B������
B���>�3���}�pz��������C��F���������=�	Y=�J��O=�C���pCOLLECT_=��+��rR���EN�/@�u�����NDE�����s#��1234567890[���!S�Y�k�F�
 %�}�)�� �߱�߷������ T��1�C��g�y�� �������,���	�� t�?�Q�c��������� ������L5֯!;2�� �9�IO  D�����v����TMRr�2!�� �	1
-��"�<����_MORz#w� ����<��� �/�%/+�m�{�$�,��?������x#+�K�$+���R�=�%�ϱ/�!�"C4/  A�&:�+�=��A{ Cz  B�� $�B�"�  �@�"�+�+�:�dڍ <#�
!5<�!99?#3�!�I=�&�-?U3z'�ݑ/Qd�!T_D[EFzA �+%J8�?�$� NUS<A���0��4KEY_TB�L  ��6��	
��� !"�#$%&'()*�+,-./d�:;�<=>?@ABC��0GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾�����A���͓��������������������������������������������������?������p�0�LCK�<��0�0S�TA��$_AUT/O_DO��&^S�IND�M^��R_3T1h_ZWT2�_����_�TRL�0L�ETE�w�Z_S�CREEN ~͚kcsc��U�MMENU ;1(�{ <o}�? |o�%[o�o�oi�o�o �o�o&�o5nE W�{����� "���X�/�A���e� w���֏�������� B��+�Q���a�s��� ������͟ߟ�>�� '�t�K�]��������� �ɯۯ(����^�5� G�m���}���ܿ��ſ ����!�Z�1�Cϐ� g�y��ϝϯ�����π��D��-�z�Q�;c_?MANUAL�_�Q�DBcjf4YDB�G_ERRL�09)Jk� ����'�9���NUML�IMc�1�%T0D�BPXWORK 1*Jk���������SDBTB_��Q +���#4��$oDB_AW�AY���GCP� �"=�S15�_A!LU�M_3���Y�Pet� ��_�� 1,�h 
���������6��_M�PISJPB��@� 	ONTIM6g��$�)��
�5��MOTNE�ND�?��RECO�RD 12Jk y����#G�O�� ��+B���!� )P�t���� Si�a/�:/L/ ^/p//�//�/'/�/ �/ ??�/6?�/Z?�/ ~?�?�?�?#?�?G?�? k? O2ODOVO�?zO�? �OO�O�O�O�OgO_ �O_�Od_v_�_�_	_ �_�_�_�_c_o*o<o �_`oKo�_�oo�o�o �ouo�o�o8�o\ n�-�%�I ��"�4��X��|�������ď֏E�3�TOLERENC@�sBȉ�N�L�����CSS_CNST_CY 23w����	ُ���A�O�a�s� ��������џߟ�� �'�9�K�a�o�������DEVICE ;24,� �� ��
��.�@�R�d�v���������HNDG�D 5,� �Cz�����LS 26ͭ���.�@�R�d��vψϮ��PARAM 7��p�՚��
��SLAVE �8ͽ��_CFG� 9�Ϛ�d�MC:\�L%0?4d.CSV�χ�cA߆�v�A n�C	Hv�߱���΁߶�
�������������<���JP��������_CRC_OUT :ͭ���_NOCOD���;����SGN� <�#M��05-JU�N-24 11:c46q�Ѯ�03q��� X�Xl���������M���Þ�j�������VERSI�ON ��V4.2.10���EFLOGIC {1=,� 	���Ё���c�PR?OG_ENBtն���ULS4 Զ�c�_ACCLIM^5��Ö��WRSTJNTT~�c�MO���ш��1INIT >�,��� /OP�T�� ?	nG
� 	R575��Û 74�	6�7R�5W��1�2�����]�~TO  ����D^�VU DKEXd('�\PATH A��A\J����H�CP_CLNTI�D ?A��� �뒃���IAG_GRP 2C�� v� 	� @K�@�G�?���?l?��>�X!* E �p/,m!���/>�.?�b�?v��"�i�^?�Vm?�Sݘ)f4�03 6789012345�"@D �� F s��@�nȴ@i�#@�d�/@_�w@�Z~�@U/@�O�@I��@�D(�*	0'�@�bn�pn�I1�A��Y�q�B4,ڠ�$�'�
21.0-�@)hs@$���@ bN@��@0���@�D@+ j
A?S?e4j
y0j	�>�R��@N@�I�@D�@�>�y@9��@�42@.v�@(��@"�\�?�?�?��?O�8L�@G�l�@BJ@<�z�@600�`�@*&@$�@�@�LO^OpO�O|�O�8=q@0��F@|�@�33@�R@�-?���?��`?�+�O��O�O_ _2\�R�@��-@&�@��@*0�!?�??� �d_v_ �_�_�_�78m`oroPo �o�o2o|o�o�o�o  &�o�on�^� �@�rE!1�15A��AMQ�P�.�� !�Y�R ��?�z�0�`-5AFH�4��N���L4Ry�X�`-@�p�p��Q�x�-r�����@�`]0Ahf'=�H�9=Ƨ�=ߺ^5=Ȯ����>�`-=��,ԏ�,�� ��'�Ca0<(�U��� 4D"Q ��-�)A@&�?h%� Z��}h�����l��� ֟p����0�B��y�>��yd��R�=���=��z�t�`-��G���G�`-p�p�aa`�Ť�@q��"@�b,�u�Bʂ `B��B��B%��`-(�/��'��V�pfb�V����\f�u!e1��c+��B��BjW�B{0AW�@���8/ݿ'�<��#�31=�4�Cw�31>
�kд�{�r�4�|���C�!����B��W��B#�Mψ8�q�$��ϒ�)� ��3����R�6��\���Xπ���%��"�[�j#������8�?���Y'ῼ�\?���}_߭�"!�CT_CONFI�G D|����eg�"!STB_F_TTS
�����8���E�m�M�AU ����MSW�_CF��E/+  �a0(�OCVIEWf�F_�k!��/ ����������� �� 4�F�X�j�|������ ����������0B Tfx��+�� ���>Pb t��'���� //(/�L/^/p/�/ �/�/5/�/�/�/ ??,$?��RCX�G�u,�!�/2>\?�?�?�?�?��?�?�?�SBL_�FAULT H�O:t�AGPMSK��*G��TDIAG� I��3�������UD1:� 6789012345�B��{A��25P���O�O�O�O__ /_A_S_e_w_�_�_�_��_�_�_�FwF29=�
��O+o��TRECP`OrJ
�Dro�G3k�O �o�o�o�o�o, >Pbt�������_oo�u�UM�P_OPTION!�#N0�TRX��'I�Q�PME �D�Y�_TEMP  _È�3B����9�����UNI=�����L�YN_BRK� J��u�EDI�TOR6�<�~��_~H`ENT 1KO9�  ,&I�RVIS:�?��{&SUMIR <���&PICK ;���&�?ʟ�������ܟ� �(� O�6�s�Z�������ͯ �����'��K�2� D���h�������ۿ¿ ���#�5��Y�@�}������EMGDI_STA��c᥁��NC_INFO �1L_���������������ì�1M_� ��9�,��
�d��ߥ߷��� �������#�5�G�Y� k�}���������� ���^�$�6�H�Z�h� ��h������������� ��0BTfx �������p� �'9K]w��� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/?1?C? U?oy?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O ?�O)_;_M_g?]_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o__!3 E�oq_{���� �����/�A�S� e�w���������я� �o�+�=�O�is� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ���#� 5�G�a�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Y�K� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������� %�7�Q�c�m������ ����������!3 EWi{���� ����/A[� ew������ �//+/=/O/a/s/ �/�/�/�/�/G�? ?'?9?S]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�/�O__1_K? U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�O�o )C_9_q� �������� %�7�I�[�m������ ��Ǐ�o�o���!�׏ MW�i�{�������ß ՟�����/�A�S� e�w���������ُ� ����+�E�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ���������#� =�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��5�'�Q�c� u��������������� );M_q� ������� -�?�I[m�� �����/!/3/ E/W/i/{/�/�/�/� ��/�/??7A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O#?�/�O�O_ _/?9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �O�o�o�o'_1C Ugy����� ��	��-�?�Q�c� u��������o���� ��;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��Ϗٯ�����)�3� E�W�i�{�������ÿ տ�����/�A�S� e�wωϛϵ�ǯ���� ���!�+�=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy������ ���-?Qc u������� //)/;/M/_/q/�/ �/��/�/�/�/	 %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�/�/�O �O�O�O?_/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�O�O�o�o�o�o_ '9K]o�� �������#� 5�G�Y�k�}����o�� ŏ׏���1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ��� ��)�;�M�_�q��� ������˿ݿ��π%�7�I�[�m�ϙ� ��$ENETMO�DE 1N���  ����������˨�R�ROR_PROG %��%���(����TABLE  ���g�yߋߙ����SEV_NUM� ��  ��������_AUT�O_ENB  ��Ž���_NO�� �O������ W *������	����+�,�>�P���FLTR����H�IS�ӧ�����_A�LM 1P�� e���죠+Q������"�4�F�U�_\����  ��������TCP_V_ER !��!��V�$EXTLOGo_REQ��������SIZ����ST�K	����T�OL  ��Dzޔ��A ��_BWDk�@ p�l��U�DIZ Q���p�ħ�qST�EP����� OP�_DO%��FDR_GRP 1R��v�d 	��#���n&���c�?��$,�MT� ��$ ���Wiz�dBkH�B��<z�������//</'/`/�A*�HkAoFa>��j/��
 E��� ��!��@R�/���/T/�/�/�?�A@� <0@�/33@�E0I3=�@@1d??�?�?F@ �5�!�!�1�>��L�FZ!D��`�D�� BT��@���{=�?�  O�?6����+B��5�?Zf5�ES;A{=����E��^*� �X���w���m�.�FE�ATURE S���l ��H�andlingT�ool �E���English �Dictiona�ry�G4D StΗ@ard�F�EAn�alog I/O��G�Ggle Sh�ift�Outo �Software UpdateY�matic Ba�ckup�IHQgr�ound Edi�t�@�GCamer�a�@F�OCnrR�ndImMS�\om�mon caliOb UIS�VnfQ��PMonitor��[tr�@Reli�ab	P�HDHCP��Y�Zata Ac�quis�S�Yia�gnosDQ�Ako�cument V�iewe�R�Wua�l Check ?Safety�Q�F?hanced�V�J��esc`FrwP�Gxt. DIO �PsfiGd�gend�`Err�PLFb�m�g%s�ir�@�` [ �J�FCTN Men�u|`v�S-wTP ;InpfacCu�E�GigEU~gu_Pp� Mask Ex�c�`g�gHTSpProxy Svdd��vigh-Spe�`Ski�T�u?`�`�mmunicCPons�xur:ppo��AVrconnecwt 2�ncrUp�stru�B
�3�e�Zat`JFe�DKAR�EL Cmd. �L�pua�xj�Ru�n-Ti�`Env�`�pel +GPs�EPS/W�GLic�ensevccl�`B�ook(Syst�em)�JMACR�Os,�r/OffseP�H�`-P
o��MR�P�REnMe�chStop�qt�#�+b�i�b[_�x��`�@EP�od
Pw�itch��3�:a.<���Optmş3�N�pfilcl2�g�~�ulti-T�p�iS�IPCM fu	n=�;�o(dwb4�[�/Regi�r�p>��ri\`FK����@N?um SelW���>�` Adju�p��x֡Z�tatu�����^j�ERDM R�obot�@sco3ve�A;�ea,��`�Freq Anl�y�wRemU��an��G;�G�Servo��`���HSNPX �b��^SNSpCl�i[a��RLibr��C޿�@ f�𰪶ozɀt:pssag4���D�� "S��K��/�IT}7�MILIB�`�:�P Firmt+RJ�P:sAcc`P�h[TPTXo8�eln�}�;��A�K��orqu
Pimu�la�Q}Q��u��PAa��J�_P�Q��&�pgev.7�#Prit`���USB po�rt �PiP�`a�\`��R EVNT�zߌ�nexcep�t�`|�i��մh�mVEC�Qr�r�r[�V'`������SѰS9C��K�SGE`�V��UI�KWeb Pl�����p�d�ZavZDT Ap�pl�t�J�֯��G�ridK�playP�G�LT)�R��.�J�c�:a ﺂ0�3Q20�0i(t�Glarm Cause/z��ed�HAscii<�qբLoadc`��gUpl���^yc	P`����uЁ`.vRA?�0�`��DZ�inAÞ���HNRTL�ϬCO}n�@e Hel�X�?�U>�����T�tr��kROS Eth��t?�$�vz���v�2D��Pkg8Upg�@ �V"�3D T�ri-_a>A��D�ef#�>Ba�d�e^����[Im�ĐF��[��nsp�#�6�64MB �DRAMo%#FR9O./tPell�L�]#sh_!k/}'c�z%�(PpA֏,ty	Ps��	b�ݐ.k{��a�R�Mmaiu`Ի�mhF����Pq+�lu��Hz�Sp�R�OzL� Sup�������0�`�pcro�F��W�x����O1uest�CrtsaF�|�L O�z���K,Pl� Bui,�n��A'PLC,OvEV�E��sCGe�OCRG�ObV�DG��O�DLS�O&V�BU_V�K��+_&Y�TAOUVB__qWp��nZi�_TCB�_��V{_�W{��W�eoT�C�O�W_�W��coTEHxo�f�O�gm�oTE_�UVF�_�g�_UVG�_1w1w[oUVHsUVIA��v�&UVLN��UMW�w�?o�wC_UVN�UVP��e�;UVRUVS������UVWߏ�S��U�VGF�)�P2 �OE��E�3�E��_D�	D��E�F#oE��D��R���TUT��0�1�)�23�)�TB�GGk�S�rain�/�UIې�HMI���pon��b����f�
"iFÌ
&�KAREL.�ݯTP_���5��"�� +�X�O�a��������� ���߿���'�T� K�]ϊρϓϥϷ��� ������#�P�G�Y� ��}ߏߡ߳������� ���L�C�U��y� �����������	� �H�?�Q�~�u����� ��������D ;Mzq���� ��
@7I vm����� /�/</3/E/r/i/ {/�/�/�/�/�/?�/ ?8?/?A?n?e?w?�? �?�?�?�?�?�?O4O +O=OjOaOsO�O�O�O �O�O�O�O_0_'_9_ f_]_o_�_�_�_�_�_ �_�_�_,o#o5oboYo ko}o�o�o�o�o�o�o �o(1^Ugy �������$� �-�Z�Q�c�u����� ������� ��)� V�M�_�q��������� �ݟ���%�R�I� [�m���������ٯ ���!�N�E�W�i� {�������޿տ�� ��J�A�S�e�wϤ� �ϭ���������� F�=�O�a�sߠߗߩ� ���������B�9� K�]�o�������� ������>�5�G�Y� k������������� ��:1CUg� ����� �	 6-?Qc��� �����/2/)/ ;/M/_/�/�/�/�/�/ �/�/�/?.?%?7?I? [?�??�?�?�?�?�? �?�?*O!O3OEOWO�O {O�O�O�O�O�O�O�O &__/_A_S_�_w_�_ �_�_�_�_�_�_"oo +o=oOo|oso�o�o�o �o�o�o�o'9 Kxo����� ����#�5�G�t� k�}���������׏� ���1�C�p�g�y� ������ܟӟ��	� �-�?�l�c�u����� ��دϯ����)� ;�h�_�q�������Կ ˿ݿ
���%�7�d��[ς�  �H552rØ�21n��R78��50���J614��ATU]P��545��6���VCAM��CRIn��UIF��28�ƷNRE��52��R�63��SCH��DwOCVR�CSU���869��0��EI�OC.�4��R69���ESET����J�7��R68��MA{SK��PRXY�]7��OCO��3��h�ƺ���3��J6���53u�H'�LCH^��OPLG��0�MHCR��Sp�MkCS��0��55���MDSW���OP��MPR�B�5�0n��PCM�R0 ������z�5�51��5u11�0��PRS�׻69��FRD��FwREQ��MCN��{93��SNBA:�^(�SHLB��M��tBЭ�2��HTC���TMIL��u�TP�A��TPTX��EL��z�u�8�ǲ���wJ95!�TUT�95��UEV��U�EC��UFR��V�CC�O��VIP���CSC!CSGt-�g�I��WEB��7HTT��R68�C�CG�IG�IP�GSRC��DG��H75��R66�Y7��R/�2�R�?��%�4��b��R�64��NVD��R6|�R84�\��6Y865�90Q�כJ9(�91)�7X ���!�D0�Fk(�CLI����CMS��֚ ��STY�T�O�7t�NN��O�RS��J��_�O]L�(END��L��S�(FVR��V3�D��PBV!A�PL��APV�C�CG��CCRq�C�D�CDL5CS�Bi�CSK��CTCTB�9��0�(�C���0�8C�TC���0u7TC�7TC���CTEQ�J@�7T�E]�J@�TF�8FJ�(G�8G�I5HH5H�I���@5H,CTM��(M)HM�8N5HP��HP�8R�8�(TSr�8WIY5VGFaWP2�P2��vPmX��7VPDmXF�V�P�GVPR6VT����P��VTB�7Vh�IH��V>�H�'VK�V�y�@oRo dovo�o�o�o�o�o�o �o*<N`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO�tO�C  H55�T|A�A�U�C�R78�L50�IJw614�IATU	d��D545�L6�IVsCAyT�CCRI![�UI�T�E28"ZN�RE�J52ZR6�3�KSCH�IDO�CV�ZC�U�D86u9�K0�JEIO!d�hU4�JR69ZEgSET�K[J7[�R68�ZMASK^�IPRXYB\7�JOCOl3�L�J`��L3qjJ6�L53��ZH�lLCHQjO�PLG�K0�jMH�CRRjS{MCS��L0!k55�JMD�SWr{�kOP�kM�PR�j~P�l0�JPCMAZR0�{`�Jlp�k51[51��0ZPRSk69�qjFRD1ZFRE�Q�JMCN�J93��JSNBAr[�kSHLB��MЋ~Pa|�2�JHTC�JTMsIL�L�ZTPA�ZoTPTX�EL���p�[8�K�@�ZJ9�5QZTUT�k95�qjUEVjUEC�QjUFR1ZVCC��O1zVIP!�C;SCQ�CSGaZ�P�I�IWEB�JHT�T�JR6p\�CG�p�IGP�IPGS���RC!�DG�kH�75ZR66�7* kR�2�jR�l�P��4qj���JR64n�ZNVDjR6 {�R84����>`�8�6�k90���[J9&�l91�A�7P[>`�QZD0p�F_�CL9I�| [CMS�Z��n�JSTY!�TOq��7�\NNqjORSb1zJ��BjO�OL��WEND�JL �S��wFVR�ZV3D!��@[PBVQ�APL��ZAPV�jCCGn�JCCRzCD �wCDL��CSB�Z�CSK�zCT@�CCTB1�Q�>���Cъ4n�1�CA�TCAZn���TC�TCjCcTE�Z����TE�Z���1�TFQ�F��GR1�G1���H��I���~���`�CTM��M���M!�N��P��P�1�RQ��TSQ�W�1��VGFQP2��P2��n ap�VkPDaFAZVP��7VPRA�VT�K� ��JVTB��V�[I�H�VΠ����VK!�Vp��Hx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O�PObOtO�C�@�STD�DLANG�D�I�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ����'�9�K�RB=T�FOPTNb�t� ��������Ο������(�:�L��EDPN �Dp���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬߀����������*� }HH�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ�������1�C�U�g�y�99�~��$FEAT_�ADD ?	��������  	}Ⱦ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4��F�X�j�|�������D�EMO S��   }��ݏ ���%�R�I�[��� ��������ٟ�� �!�N�E�W���{��� ����ޯկ���� J�A�S���w������� ڿѿ����F�=� O�|�sυϟϩ����� �����B�9�K�x� o߁ߛߥ�������� ���>�5�G�t�k�}� ������������� :�1�C�p�g�y����� ������ ��	6- ?lcu���� ���2);h _q������ �/./%/7/d/[/m/ �/�/�/�/�/�/�/�/ *?!?3?`?W?i?�?�? �?�?�?�?�?�?&OO /O\OSOeOO�O�O�O �O�O�O�O"__+_X_ O_a_{_�_�_�_�_�_ �_�_oo'oToKo]o wo�o�o�o�o�o�o�o #PGYs} �������� �L�C�U�o�y����� ��܏ӏ��	��H� ?�Q�k�u�������؟ ϟ����D�;�M� g�q�������ԯ˯ݯ 
���@�7�I�c�m� ������пǿٿ��� �<�3�E�_�iϖύ� ������������8� /�A�[�eߒ߉ߛ��� ���������4�+�=� W�a��������� �����0�'�9�S�]� ���������������� ��,#5OY�} �������( 1KU�y�� �����$//-/ G/Q/~/u/�/�/�/�/ �/�/�/ ??)?C?M? z?q?�?�?�?�?�?�? �?OO%O?OIOvOmO O�O�O�O�O�O�O_ _!_;_E_r_i_{_�_ �_�_�_�_�_ooo 7oAonoeowo�o�o�o �o�o�o3= jas����� ����/�9�f�]� o�������ҏɏۏ� ���+�5�b�Y�k��� ����Οşן���� '�1�^�U�g������� ʯ��ӯ ���	�#�-� Z�Q�c�������ƿ�� Ͽ�����)�V�M� _όσϕ��Ϲ����� ����%�R�I�[߈� ߑ߾ߵ��������� �!�N�E�W��{�� ������������� J�A�S���w������� ��������F= O|s����� ��B9Kx o������� //>/5/G/t/k/}/ �/�/�/�/�/�/?? :?1?C?p?g?y?�?�? �?�?�?�?�?	O6O-O ?OlOcOuO�O�O�O�O �O�O�O_2_)_;_h_ __q_�_�_�_�_�_�_ �_o.o%o7odo[omo �o�o�o�o�o�o�o�o *!3`Wi�� ������&�� /�\�S�e�������ȏ ��я���"��+�X� O�a�������ğ��͟ ����'�T�K�]� ����������ɯ�� ��#�P�G�Y���}� ������ſ߿��� �L�C�Uς�yϋϸ� ���������	��H� ?�Q�~�u߇ߴ߽߫� �������D�;�M� z�q��������� 
���@�7�I�v�m� ������������� <3Eri{�|��  � ��);M_ q������� //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o����������ɉ  ʈρ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w�����(����΁Ӏƈ� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew�����	�$FE�AT_DEMOIoN  ����� �INDE�X��� IL�ECOMP T����7��-SETUPo2 U7A?�  N l*�_AP2BCK �1V7  �)���%��� :����*/� N/�[/�//�/7/�/ �/m/?�/&?8?�/\? �/�?�?!?�?E?�?i? �?O�?4O�?XOjO�? �OO�O�OSO�OwO_ _�OB_�Of_�Os_�_ +_�_O_�_�_�_o�_ >oPo�_too�o�o9o �o]o�o�o�o(�oL �op��5�� k ��$�6��Z�� ~������C�؏g��� ���2���V�h����� ���Q��u�
��� �@�ϟd�󟈯��)� ��M���������<� N�ݯr����%���̿tFzP~ 2�*.VRӿϋ�* �Fψ�L�p�Z���PCxϡϋ�F'R6:����\�����T�'߶��Q��� ��w�Y�*.F�
Ϩߊ�	�Ö���8d��߈�STM�.��»��Y���}��HJ��?��[�m����GIF�6�A�"�p�������JPG�����A��c�u�
��JS=����+���%
JavaSc�ripti��CS�Z�@�k %�Cascadin�g Style ?Sheets�_��
ARGNAME�.DT�D�\@0�P`q`DISP*gJD��������
T�PEINS.XML$/�:\8/�X�Custom T?oolbary/��PASSWORD��}�FRS:\��/{/ %Pas�sword Config�/X�F?�/ ??|?���?/?�?�?e? �?�?O0O�?TO�?xO OO�O=O�OaO�O_ �O,_�OP_b_�O�__ �_�_K_�_o_o�_�_ :o�_^o�_Wo�o#o�o Go�o�o}o�o6H �ol�o�1�U �y� ��D��h� z�	���-�ԏc��� �������R��v�� o���;�П_������ *���N�`����� 7�I�ޯm������8� ǯ\�므���!���E� ڿ�{�ϟ�4�ÿտ j�����χ���S��� w��߭�B���f�x� ߜ�+���O�a��߅� ���P���t��� ��9���]������(� ��L���������5� ����k� ��$6�� Z��~��C� gy�2�+h ����Q�u 
//�@/�d/�/ �/)/�/M/�/�/�/? �/<?N?�/r??�?�? 7?�?[?�??�?&O�? JO�?CO�OO�O3O�O �OiO�O�O"_4_�OX_��O|___�_�V�$�FILE_DGB�CK 1V����P��� < �)
SU�MMARY.DG<�_h\MD:�_0o�tPDiag Summary1o�>Z
CONSLO�G&o	oato�oCa�Console �log�o=[	TPOACCN�o%�o�4?eTP Accountin�o�>ZFR6:IP�KDMP.ZIP�hlX
��@ePpE�xception��n{`MEMCH�ECK*�oo@���aMemory �DataA��V-�l�)+�RIPE�o�+���O�%��� Packet� L�o�TL�$�<�r��STAT����|��H� %܂?StatusI���	FTP����/����K��amment� TBD͟�� >�I)ETHERNE����q�P�CaEthern�~�`figura��DT��DCSVRF�������үY��� �verify a�llկ�SM.���DIFFʯ��¯xW�փ�diffY����q��CHG01 N�5�G�ܿ[�o���-?��2ҿ��˿`�k��ϡ�3V�=�Oώ�� v�ߚ��VTRNDIAG.LS�����h�S�=(� Opex��� Hanostic�u���)VD;EV,�DATi�F�xX�j�\�Vis��?Device�ߟ�IMG,ү����n�zՃ�Imag�n��UP��ES��~I�FRS:\�����DaUpdates List���>Z\�FLEXEVENF�M�_�x�[��;� UIF E�v�菖R,�s��)
PSRBWLOD.CM��h\��������`PS_RO�BOWEL�:GIG��Wb�{N�GigE����R�N�? )lHADOWv[m�Q�Shadow Changej��w�b�RCMERR����Q��KCFG Er�ror
�tail�) MA��C?MSGLIB~e�w/��d��ic����)�Z�DGf/��/M�ZMD� ad,/��NOTI��i/{/?�O�Notifiqcy��/���AGJ_ g?n_�?�_�?�?D_�? t?	OO�??O�?cOuO O�O(O�O�O^O�O�O _�O$_M_�Oq_ _�_ �_6_�_Z_�_o�_%o �_Io[o�_oo�o2o �o�oho�o�o!3�o W�o{��@� �v��/��<�e� ��������N��r� ����=�̏a�s�� ��&���J�ȟ񟀟� ��9�K�ڟo������� 4�ɯX������#��� G�֯T�}����0�ſ ׿f������1���U� �yϋ�ϯ�>���b� ��	ߘ�-߼�Q�c��� ��߽߫�L���p�� ��;���_���l�� $��H�����~���� 7�I���m������2� ��V���z���!��E ��i{
�.�� d��/�S� w��<�`� /�+/�O/a/��/ /�/�/J/�/n/?�/ ?9?�/]?�/�?�?"? �?F?�?�?|?O�?5O GO�?kO�?�OO�O�O��C�$FILE_�FRSPRT  ����@�����HMDO?NLY 1V�E�@� 
 �)�MD:_VDAEXTP.ZZZ�O�}OT_c[6%�NO Back �file ._�DS�6PZO�_D_�_�O �_oTO3o�_Woio�_ �oo�o�oRo�ovo �oA�oe�or� *�N����� =�O��s������8� ͏\�񏀏��'���K� ڏo������4�ɟ۟�j�����#�5��DVI�SBCKX�AS�*.VD6�����FR:\O�ION?\DATA\k����Vision VD�R������ ��*��N�ݯ_��� ���7�̿޿m�ϑ� &ϵ�ǿ\�뿀ϒ�M� ��E���i���ߟ�4� ��X�j��ώ�߲�A� S���w�����B��� f���w��+���O��� ������>�����t���JLUI_CON�FIG W�E�b�� $  ]��C������ $<6T$ |xf�h z����V�� +�<as� ��@���// '/�K/]/o/�/�/�/ </�/�/�/�/?#?�/ G?Y?k?}?�?�?8?�? �?�?�?OO�?COUO gOyO�O�O4O�O�O�O �O	__�O?_Q_c_u_ �__�_�_�_�_�_o �_)o;oMo_oqo�oo �o�o�o�o�o�o% 7I[m�� �����!�3�E� W�i�{������ÏՏ ������/�A�S�e� w��������џ�z� ���+�=�O�a����� ������ͯ߯v��� '�9�K�]��������� ��ɿۿr����#�5� G�Y��}Ϗϡϳ��� ��n�����1�C�U� ��yߋߝ߯�����j� ��	��-�?���P�u� �����T������ �)�;���_�q����� ����P�����% 7��[m��� L���!3� Wi{���D����////� � x;/H#�$F�LUI_DATA X���x!��j$R�ESULT 2Y�x%�  �T��W/�/�/�/�/? ?)?;?M?_?q?�?�? ��/�?�?�?�?OO )O;OMO_OqO�O�O�O��M?�0��x%�O�K��_"_ 4_F_X_j_|_�_�_�_ �_�_�_�3�Oo$o6o HoZolo~o�o�o�o�o�o�o�{ �Ow�O 0�OWi{��� ������/�A� Re�w���������я �����+�=��o^�  ��D����͟ߟ� ��'�9�K�]�o��� ��R���ɯۯ���� #�5�G�Y�k�}���N� ��r�Կ������1� C�U�g�yϋϝϯ��� ���Ϥ�	��-�?�Q� c�u߇ߙ߽߫����� ���Ŀ&�8���_�q� ������������ �%�7���[�m���� ������������! 3��<��`�L� ����/A Sew�H���� ��//+/=/O/a/ s/�/D�h�/�/� ??'?9?K?]?o?�? �?�?�?�?�?��?O #O5OGOYOkO}O�O�O �O�O�O�/�/�/�/._ �/U_g_y_�_�_�_�_ �_�_�_	oo-o�?Qo couo�o�o�o�o�o�o �o);�O__ �B_������ �%�7�I�[�m��>o ����Ǐُ����!� 3�E�W�i�{���L^ pҟ�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿��  �$��K�]�oρ� �ϥϷ���������� #�5�F�Y�k�}ߏߡ� ������������1� �R��v�8ϝ���� ������	��-�?�Q� c�u���F߫������� ��);M_q �B�f���� %7I[m� �������/!/ 3/E/W/i/{/�/�/�/ �/�/��/�?,?� S?e?w?�?�?�?�?�? �?�?OO+O�OOaO sO�O�O�O�O�O�O�O __'_�/0?
?T_~_ @?�_�_�_�_�_�_o #o5oGoYoko}o<O�o �o�o�o�o�o1 CUgy8_�_\_� ��_�	��-�?�Q� c�u���������Ϗ�o ���)�;�M�_�q� ��������˟��� �"��I�[�m���� ����ǯٯ����!� ��E�W�i�{������� ÿտ�����/��  ��t�6��ϭϿ��� ������+�=�O�a� s�2��ߩ߻������� ��'�9�K�]�o�� @�R�d��������� #�5�G�Y�k�}����� ����������1 CUgy���� ��������?Q cu������ �//)/:M/_/q/ �/�/�/�/�/�/�/? ?%?�F?j?,�? �?�?�?�?�?�?O!O 3OEOWOiO{O:/�O�O �O�O�O�O__/_A_ S_e_w_6?�_Z?�_~? �_�_oo+o=oOoao so�o�o�o�o�o�O�o '9K]o� �����_��_�  ��oG�Y�k�}����� ��ŏ׏������o C�U�g�y��������� ӟ���	���$�� H�r�4�������ϯ� ���)�;�M�_�q� 0�������˿ݿ�� �%�7�I�[�m�,�v� P����φ������!� 3�E�W�i�{ߍߟ߱� �߂�������/�A� S�e�w�����~� �Ϣϴ����=�O�a� s��������������� ��9K]o� ������� #�����h*��� �����//1/ C/U/g/&�/�/�/�/ �/�/�/	??-???Q? c?u?4FX�?|�? �?OO)O;OMO_OqO �O�O�O�Ox/�O�O_ _%_7_I_[_m__�_ �_�_�_�?�_�?o�? 3oEoWoio{o�o�o�o �o�o�o�o.oA Sew����� �����_:��_^�  o��������͏ߏ� ��'�9�K�]�o�. ������ɟ۟���� #�5�G�Y�k�*���N� ��r�t������1� C�U�g�y��������� �����	��-�?�Q� c�uχϙϫϽ�|��� ����ؿ;�M�_�q� �ߕߧ߹�������� �ҿ7�I�[�m��� �������������� ���<�f�(ߍ����� ��������/A Se$����� ��+=Oa  �j�D���z��� //'/9/K/]/o/�/ �/�/�/v�/�/�/? #?5?G?Y?k?}?�?�? �?r���
O�1O COUOgOyO�O�O�O�O �O�O�O	_�/-_?_Q_ c_u_�_�_�_�_�_�_ �_oo�?�?�?\oO �o�o�o�o�o�o�o %7I[_� �������!� 3�E�W�i�(o:oLo�� poՏ�����/�A� S�e�w�������l�� �����+�=�O�a� s���������z�ܯ��  �'�9�K�]�o��� ������ɿۿ���� "�5�G�Y�k�}Ϗϡ� �����������̯.� �R��yߋߝ߯��� ������	��-�?�Q� c�"χ�������� ����)�;�M�_�� ��Bߤ�f�h����� %7I[m� ��t����! 3EWi{��� p�����/�//A/ S/e/w/�/�/�/�/�/ �/�/?�+?=?O?a? s?�?�?�?�?�?�?�? O�/�0OZO/�O �O�O�O�O�O�O�O_ #_5_G_Y_?}_�_�_ �_�_�_�_�_oo1o CoUoO^O8O�o�onO �o�o�o	-?Q cu���j_�� ���)�;�M�_�q� ������foxo�o�o�� �o%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ����ʏ܏� P��w���������ѿ �����+�=�O�� sυϗϩϻ������� ��'�9�K�]��.� @���d���������� #�5�G�Y�k�}��� `ϲ���������1� C�U�g�y�������n� ��������-?Q cu������ �);M_q �������/ ��"/��F/m//�/ �/�/�/�/�/�/?!? 3?E?W?{?�?�?�? �?�?�?�?OO/OAO SO/tO6/�OZ/\O�O �O�O__+_=_O_a_ s_�_�_�_h?�_�_�_ oo'o9oKo]ooo�o �o�odO�o�O�o�o�_ #5GYk}�� ������_�1� C�U�g�y��������� ӏ����o �o$�N� u���������ϟ� ���)�;�M��q� ��������˯ݯ�� �%�7�I��R�,�v� ��b�ǿٿ����!� 3�E�W�i�{ύϟ�^� ����������/�A� S�e�w߉ߛ�Z�l�~� ���ߴ��+�=�O�a� s����������� ���'�9�K�]�o��� ���������������� ����D�k}�� �����1 C�gy���� ���	//-/?/Q/ "4�/X�/�/�/ �/??)?;?M?_?q? �?�?T�?�?�?�?O O%O7OIO[OmOO�O �Ob/�O�/�O�/_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_
_o/oAo Soeowo�o�o�o�o�o �o�o�O�O:�Oa s������� ��'�9�K�
oo��� ������ɏۏ���� #�5�G�h�*��N P�şן�����1� C�U�g�y�����\��� ӯ���	��-�?�Q� c�u�����X���|�޿ 𿴯�)�;�M�_�q� �ϕϧϹ������Ϯ� �%�7�I�[�m�ߑ� �ߵ������ߪ���ο �B��i�{���� ����������/�A�  �e�w����������� ����+=��F�  �j�V���� '9K]o� �R������/ #/5/G/Y/k/}/�/N `r��/�??1? C?U?g?y?�?�?�?�? �?�?�	OO-O?OQO cOuO�O�O�O�O�O�O �O�/�/�/8_�/__q_ �_�_�_�_�_�_�_o o%o7o�?[omoo�o �o�o�o�o�o�o! 3E__(_�L_� ������/�A� S�e�w���Ho����я �����+�=�O�a� s�����V��zܟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿鿨�
�̟.� �U�g�yϋϝϯ��� ������	��-�?��� c�u߇ߙ߽߫����� ����)�;���\�� ��B�D��������� �%�7�I�[�m���� Pߵ���������! 3EWi{�L� p�����/A Sew����� ���//+/=/O/a/ s/�/�/�/�/�/�/� ��?6?�]?o?�? �?�?�?�?�?�?�?O #O5O�YOkO}O�O�O �O�O�O�O�O__1_ �/:??^_�_J?�_�_ �_�_�_	oo-o?oQo couo�oFO�o�o�o�o �o);M_q �B_T_f_x_��_� �%�7�I�[�m���� ����Ǐُ�o���!� 3�E�W�i�{������� ß՟矦��,�� S�e�w���������ѯ �����+��O�a� s���������Ϳ߿� ��'�9���
��~� @��Ϸ���������� #�5�G�Y�k�}�<��� ������������1� C�U�g�y��JϬ�n� �����	��-�?�Q� c�u������������� ��);M_q ��������� ��"��I[m� ������/!/ 3/��W/i/{/�/�/�/ �/�/�/�/??/?� P?t?68?�?�?�? �?�?OO+O=OOOaO sO�OD/�O�O�O�O�O __'_9_K_]_o_�_ @?�_d?�_�_�O�_o #o5oGoYoko}o�o�o �o�o�o�O�o1 CUgy���� ��_�_�_ �*��_Q� c�u���������Ϗ� ���)��oM�_�q� ��������˟ݟ�� �%��.��R�|�>� ����ǯٯ����!� 3�E�W�i�{�:����� ÿտ�����/�A� S�e�w�6�H�Z�l��� ������+�=�O�a� s߅ߗߩ߻��ߌ��� ��'�9�K�]�o�� ��������ϬϾ�  ���G�Y�k�}����� ������������ CUgy���� ���	-���� �r4������ �//)/;/M/_/q/ 0�/�/�/�/�/�/? ?%?7?I?[?m??> �?b�?��?�?O!O 3OEOWOiO{O�O�O�O �O�O�?�O__/_A_ S_e_w_�_�_�_�_�_ �?�_�?o�?=oOoao so�o�o�o�o�o�o�o '�OK]o� �������� #��_D�oh�*o,��� ��ŏ׏�����1� C�U�g�y�8������ ӟ���	��-�?�Q� c�u�4���X���̯�� ���)�;�M�_�q� ��������˿���� �%�7�I�[�m�ϑ� �ϵ��φ�Я����� �E�W�i�{ߍߟ߱� ����������ܿA� S�e�w������� ��������"���F� p�2ߗ����������� '9K]o.� ������� #5GYk*�<�N� `������//1/ C/U/g/y/�/�/�/�/ ��/�/	??-???Q? c?u?�?�?�?�?�?� ��O�;OMO_OqO �O�O�O�O�O�O�O_ _�/7_I_[_m__�_ �_�_�_�_�_�_o!o �?�?Ofo(O�o�o�o �o�o�o�o/A Se$_v���� ����+�=�O�a� s�2o��Vo��zoߏ� ��'�9�K�]�o��� ������ɟڏ���� #�5�G�Y�k�}����� ��ů��毨�
�̏1� C�U�g�y��������� ӿ���	��ڟ?�Q� c�uχϙϫϽ����� ����֯8���\��  ߕߧ߹�������� �%�7�I�[�m�,ϑ� ������������!� 3�E�W�i�(ߊ�L߮� ��������/A Sew����~� ��+=Oa s����z����� �/��9/K/]/o/�/ �/�/�/�/�/�/�/? �5?G?Y?k?}?�?�? �?�?�?�?�?O�/ �:OdO&/�O�O�O�O �O�O�O	__-_?_Q_ c_"?�_�_�_�_�_�_ �_oo)o;oMo_oO 0OBOTO�oxO�o�o %7I[m� ��t_����!� 3�E�W�i�{������� Ï�o�o�o��o/�A� S�e�w���������џ �����+�=�O�a� s���������ͯ߯� ��ԏ���Z���� ������ɿۿ���� #�5�G�Y��jϏϡ� ������������1� C�U�g�&���J���n� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� ��������x������� ��%7I[m� �������� 3EWi{��� ����/��,/�� P//�/�/�/�/�/ �/�/??+?=?O?a?  �?�?�?�?�?�?�? OO'O9OKO]O/~O @/�O�Ox?�O�O�O_ #_5_G_Y_k_}_�_�_ �_r?�_�_�_oo1o CoUogoyo�o�o�onO �O�O�o�O-?Q cu������ ���_)�;�M�_�q� ��������ˏݏ�� �o
�o.�X���� ����ǟٟ����!� 3�E�W��{������� ïկ�����/�A� S��$�6�H���l�ѿ �����+�=�O�a� sυϗϩ�h������� ��'�9�K�]�o߁� �ߥ߷�v������߾� #�5�G�Y�k�}��� ������������1� C�U�g�y��������� ������	������N �u������ �);M�^ �������/ /%/7/I/[/|/> �/b�/�/�/�/?!? 3?E?W?i?{?�?�?�? �/�?�?�?OO/OAO SOeOwO�O�O�Ol/�O �/�O�/_+_=_O_a_ s_�_�_�_�_�_�_�_ o�?'o9oKo]ooo�o �o�o�o�o�o�o�o�O  �OD_}�� �������1� C�U�oy��������� ӏ���	��-�?�Q� r�4����l�ϟ� ���)�;�M�_�q� ������f�˯ݯ�� �%�7�I�[�m���� ��b�����п����!� 3�E�W�i�{ύϟϱ� �������ϸ��/�A� S�e�w߉ߛ߭߿��� ���ߴ���ؿ"�L�� s����������� ��'�9�K�
�o��� �������������� #5G��*�<� `�����1 CUgy��\�� ���	//-/?/Q/ c/u/�/�/�/j|� �/�?)?;?M?_?q? �?�?�?�?�?�?�?� O%O7OIO[OmOO�O �O�O�O�O�O�O�/�/ �/B_?i_{_�_�_�_ �_�_�_�_oo/oAo  ORowo�o�o�o�o�o �o�o+=O_ p2_�V_���� ��'�9�K�]�o��� �����ɏۏ���� #�5�G�Y�k�}����� `�柨��1� C�U�g�y��������� ӯ������-�?�Q� c�u���������Ͽ� 󿲟�֟8�����q� �ϕϧϹ�������� �%�7�I��m�ߑ� �ߵ����������!� 3�E��f�(ϊ��`� ����������/�A� S�e�w�����Z߿��� ����+=Oa s��V��z��� ��'9K]o� ��������/ #/5/G/Y/k/}/�/�/ �/�/�/�/���? @?g?y?�?�?�?�? �?�?�?	OO-O?O� cOuO�O�O�O�O�O�O �O__)_;_�/?? 0?�_T?�_�_�_�_o o%o7oIo[omoo�o PO�o�o�o�o�o! 3EWi{��^_ p_�_��_��/�A� S�e�w���������я ㏢o��+�=�O�a� s���������͟ߟ� ���6��]�o��� ������ɯۯ���� #�5��F�k�}����� ��ſ׿�����1��C��d�&��ϖ��$�FMR2_GRP� 1Z���� �C4 w B�O�	 O��������F@ ��E�����H�����L�FZ!D��`�D�� BT��@���ݏ?�  L�H���6����t���5�Zf5�ES�ў�A�  �߮�B�H�����@�33K@�����H��������@������U���<�z�<��ڔ=7�<��
;;�*�<����8ۧ�9�k'V8��8����7ג	8(��4��X���������;�M���_C_FG [��T���w�������O�NO {��
F0��� ��L�RM_CHKTYP  ���O�����w���ROM���_MIN O����. ���X��S�SB]�\�� ��[O�R�{�S�TP_DEF_OW  O���âIRCOM� ��$GENO�VRD_DO#�Y��THR# dz�d�_ENB�{ � RAVC��u]DO  ��� �~,�����n�� �FOU��c�����ȷ��<+ ^�8/�0/�R/�/O�C�  D � �/"&�/�,@���,B����"��#)�GSMT��dT��Q ��$�$HOSTC�]�1e��P �\Y��� MCO��+�{?O�  2�7.0�01�?  e�?�?
OO.O<J �?_OqO�O�O�<OOIC�	anonymous�O�O�O_ _2_ z?��GXG[�?�O �_�?�_�_�_�_oKO (o:oLo^o�_o�O�o �o�o�o�o5_�oY_k_ Ho�__���� o��� �2�U�o �oz�������	 -?A�.�uR�d�v� �������П���� )�_� �N�`�r����� ݏ��ޯ��I�&� 8�J�\����������� ȿ�m�3��"�4�F� Xϟ���ïկ׿��� ������0�w�T�f� xߊߜ߿�������� ��,�sυϗ�t�� ���ϼ�������߯� (�:�L�^�����ߦ� ��������5�G�Y�k� m�?��~���� ��� 2U�� ��z����/4]1�ENT 1f+� P!K	/  +0�4/#/X//|/ ?/�/c/�/�/�/�/�/ ?�/B??f?)?�?M? _?�?�?�?�?O�?,O �?ObO%O�OIO�OmO �O�O�O_�O(_�OL_ _p_3_|_W_�_�_�_ �_�_o�_6o�_Zoo�/o�oSo�owo�o�j?QUICC0�o�o�o4�d15#���d2�as�!?ROUTER����$�!PCJO�G%� �!19�2.168.0.�10�o�cCAMP�RTu�Q�!e�1n�����RT������� !Soft�ware Ope�rator Pa�nel��b�c��N�AME !�!�ROBO��k�S_CFG 1e�� �A�uto-star�tedFTP'��>@'�tK� ]�o��������ɯۯ ������5�G�Y�k� }���՟���ֿ�/� ��0�B�T��xϊ� �Ϯ����e����� ,�>�P�);�� ���������(��� L�^�p����9��� ���� ��$�k�}ߏ� l�����ߴ������� �� 2DVy��� u�����-�?� Q�c�eR��v�� �����//*/ M�`/r/�/�/�/�/ %?9/&?mJ? \?n?�?G/=?�?�?�? �??O�?4OFOXOjO |O�/�/�/�/�?�O/? __0_B_T_Ox_�_ �_�_�_�Oe_�_oo ,o>oPo�O�O�Oio�_ �o_�o�o(�_ L^p��o�9���� ����z�_ERR g��"�2��PDUSIZ  ��p^�`�I�>~b�WRD ?Õ��a�  guest�v�����Ə؏���s�SCD�_GROUP 3�hÜ Ǒ�yI�FTB�$PAB�O�MPB� B�_�SHB�ED�� $�CB�COM4�TT�P_AUTH 1�iA� <!i?Pendan�����Ʒ!KARE�L:*��.�K�CC�S�e�;�VI�SION SET�,�ï��4�گȯ� �:��#�p�G�Y�{��}������CTRL� jA����q
���FFF9�E3���dFRS�:DEFAULT�!�FANUC� Web Server!����┊� ��ʼ�ϩϻ��������0�WR_CONF�IG k1��}�!�2�IDL_CPU_PC@���qBȕ`c� BHI�MINT�9�g�?GNR_IO;�p���pG�K�NPT_S_IM_DO�����STAL_SCR�N�� �����TPMODNTOL����|�RTY��cѨ�\���ENB��9��H�OLNK 1lA�>�k�}���������O�MASTE��?��OSLA�VE mA��RAMCACHE�����O�O_CFG7�N�O�UO Z�K�?CMT_OP@���E���YCL6�i�:�_ASG 1n&�|�
 ����  2DVhz�����������NUMjo�E�
K�IP4��F�RTRY_CNx��i���_UPDo��j��I� K�v�T��o�6��6�K�P_�MEMBERS �2p&�� $1�����S��K�RC�A_ACC 2q�1�  XŇ[����r6�M"�`�pq�A&R#L#�V/H!m/߱%"BUF001 2r1��= �gu0 _ u0�w�$��$U��$��$��$��$���$��#�4�4(484K4[�4c q� �`V�#�oD4�D4�D4U�D4�D4�D4�D4��D4��#�4���4&�45�4G�4V̌4�$�x�4�$����4�$���4ь4㬌4�4�DD)�D:DLD]Dp�D�D�D�D��D�D�D�D���$�$!�$1�$C�$T�#�)2�/�#�! �!�B� �B� �B� �B � �B� �B� �B0�! 
1R0R0R#0R +0R30R;0<1B1�! J1ORS0OR[0ORc0OR k0ORs0OR{0OR�0OR �0�!�1�R�0�R�0�R �0�R�0�R�0�R�D�1 �R�D�1�R�D�1�R�0 �R�0�R�T
Ab@b @b#@b+@b3@b ;@bC@bK@bS@b [@bc@bk@bs@b {@�B�@�B�@�B�@�B �@�B�@�!�)3�O�% �C�b�"�C�b�"�C�b �"S�b2Sr2!S r#21Sr32AS�qB3 QSPrS2aSPrc2qSPr s2�SPr�2�S�q�3�S �r�2�S�r�2�S�r�d �3�S�r�2�S�r�2�S �r�2	c��
Cc�B )c�+B9c�;BIc� KBYc�[Bic�kByc �{B�c�b�B�c�b�B��cG�&!U�2s1�C 4��Ś��!<�$p������#$HIS�"�u1� �A! �2024-06-05��i�Z�l�~�z��`֑; h�� p��x֑��l"���[��ӟ������ �G�4�F�X�j�|��� ����į֯���� 0�B�T�f�x������� ��������,�>� P�b�tφϽ�Ͽ���� ������(�:�L�^� �ϧϹϦ߸�������  ��$�6�H�ߑ�~� �������������  ���@�/�A�w������������d���� d������t ��ː ���	U�g�Qc u������� *<);M_q� ����&/ %/7/I/[/m//�/�/ �/���/�/?!?3? E?W?i?{?�?�/�/�? �?�?�?OO/OAOSO eO�?�?�O�O�O�O�O �O__+_=_+��bB� T�f��_�_�_�_���� ���R���R���RÐ �R���Ro.o@ozO�O vo�o�o�o�o�o�o�o OoaoN`r� ������'9 K8�J�\�n������� ��ȏڏ�#��"�4� F�X�j�|�������� �������0�B�T� f�x�����ӟ��ү� ����,�>�P�b�P\�I_CFG 2v�h[ H
Cy�cle Time���Busy���Idl����mi�nk�ݱUp|����Read���DowѸͿ ����Coun}t��	Num ��"�����N̉P%�3�oPROG��whUrP�^ϣϵ����������ع.�SDT�_ISOLC  �hY� =�n�J�23_DSP_ENB  0�ްQ�?INC xa݉S�>�A   ?��=���<#�
=�>��:�o �Ѽ�`�߉Q����J�OBy��CZ�ٵ���G_�GROUP 1yv0���<��P�ә�\���?������PQ��������� �0�B�T�������G_IN_AUT�O�e�POSRE��*�KANJI_�MASK������R�ELMON zh[VωRy�2DV�hzn���}�{���lӉT���m�KCwL_L��NUM^���$KEYLOGOGING� mP�P��i�t�LANGUA_GE hU8��DEFAUgLT FVQLG���|��ݲ�d���P8ްH  �V�P'0����P;�PxmಉU;��
�(UT1:\�� ���//�+/=/O/f/s/�/�.(�!�/QVLN_DISP }{�ڸ��|���$OCTOL'0��QDzn�9є�=1GBOOK ~W�d�$౨!�!u0X ��?�?�?�?�?�;M0c޳I�6	[5��X��]Oߎ�Y2_B�UFF 20� ���P2ٵ�Ot2 ��O׷�O�O__$_ Q_H_Z_�_~_�_�_�_ �_�_�_oo oMon�~�ADCS ��� �Ҝ�LQO�����o�o��o�oddIO 2��pk ��!X��$4FXl|� �������� 0�D�T�f�x����������ԏ�eER_ITM-�dr�-�?�Q�c� u���������ϟ�� ��)�;�M�_�q���8��77�SEV� a�]��TYP-������!�����RST��beSCRN_F�L 2�}n�� �o������˿ݿ��F2�TP-��1=NGNAMZԎ58n`dUPS� GIJ���i�p�_LO{AD�G %.�%SUMIR���MAXUALR�M���1@�i�
���v�_PR{ļ� hO3A��C� �e=�/��O�u1�6�P �2�e; ؟&	 쯚߅߾ߩ������� ��<��1�r�]�� ������������� 	�J�5�n�Y������� ����������"F 1j|_���� ���	BT7 xc����� �/,//P/;/t/W/ i/�/�/�/�/�/?�/ (??L?/?A?�?m?�? �?�?�?�? O�?$O���DBGDEF � Չa,�<D_LDXDISA[�-��cMEMO_APU��E ?.�
 RAH�O�O�O�O�O�__,_��FRQ_�CFG � �6VCA G@�sS@<�dd%/\�_@_RP�h҈ �D�*�P/�R **:�RD�_�X�_F o,oYoPobo�o�o�o �oO ��o��o'w,(�ol�dZ �~������ �9�K�2�o�V��������ɏ��ISC 1�.��P �O�D WO'�O`�K���Տ��_MSTR ������SCD 1��M�|���x���>� )�b�M�_��������� �˯���:�%�^� I���m�����ʿ��ǿ  ��$��H�3�l�W� |Ϣύ��ϱ������ ��2��/�h�Sߌ�w� �ߛ��߿���
���.� �R�=�v�a���� ���������<�'� L�r�]����������������MKUQ�����Q$MLTA[RMTR��W? 0sP@~�?@�METPUy@�������NDSP_ADCOL�T@�oCMNT� ��FN� ��FST�LI��� ����Uu�Qmw�P�OSCF#�PgRPM��ST� �1��� 4R#�
����/'� //#/e/G/Y/�/}/ �/�/�/�/?�/�/=?�?1?s?]1�SIN�G_CHK  �$MODASS��=?�5DEV� 	|J	MC}:�<HSIZEyM���ȭ5TASK �%|J%$123456789 NO�`E�7TRIG 1��� l?E�_�O`6y�O�O6}0FYPA�6u�4�3EM_I�NF 1��[�`)AT&FVg0E0�OY])AQ�E0V1&A3&�B1&D2&S0�&C1S0=H])�ATZY_�_�TH@�_�_hQ�Oo�XA	o@1o�_Uo<oyo�o ?_ �oc_u_�_�_
�_. eoRdo�C�� ���o�o��o�o�o `�k%�����u� �������8�J��n� !�3�E�W�ȟ{��#� ��"�ՏF��j�|�c� ��S�e�֯������� 0��T���x�3�=��� i�ҿ����ϻ�,�߯ �����9��ϼ�� �ϓ�߿��:�!�^߾�?NITOR>G� ?�;   	?EXEC1���U2��3��4��5��Tq@��7��8��9����(������ ������������@��������2�U2�2+�27�2C�U2O�2[�2g�2s�U2�3�3�3����1R_GRP_S�V 1�.[ (�e1�C��?����� � �\���?C���=8A_D��Ng�ION_DB�0�|�=��  ���8��&����q ��8T�N   �#ߵ�\�9-ud1E/A��PL_NAME �!?Ej �!�Default �Personal�ity (fro�m FD)��R�R2%� 1�L?�XL�pj�� dh��� ��#5GYk }�������//1/�32�\/n/ �/�/�/�/�/�/�/�/�2<K/(?:?L?^?p? �?�?�?�?�?�?�?I%6?(N
OLOKP;OxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_UOgO�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�_�_  $6HZl~� ������� �� H�6 H?�b H\�KA��  �M�_�Kd I�1�~���t�����2� %�H
������+�.� �F�<�N�`� ~�����ğA�����K�	`0�*�<�|N��:�oA��n������� A�  ���گ� ����1��U�g�R�Ћ�v���NR$� 1�b	���@ �� T�j � 3@D[���?����?K �KA��6�Ez  "�	4�;��	l�	 ��@�� 0<� O� ����� � �� �t�A�J���K ��J˷��J� �J�4�JR�<�������^���A�@�S�@��;fA6A���A1UA狠X�ϸ��=��N��f������T;f���X��ڮ��*�  ��  �O5��>@�[��?����?+�?��w�#�K��������ߔ������-��1ϻ�җЄ����(  ���������֢���	'�� � 2�I�� �  ��ƥ��:�ÈV�ß�=���n��߶� <O��� � � �������������� � � '����@!�p@�a�@#е@'�@+�C?�C�P��P�K�B��CzS����@���  �=ɚ�00�ɹ��i�i���@K ��KD '�� ��$H3���s���� :�Η  ��x?��ffя��X !����8��#1>�צ������^Ph�	e�^�^Ğ��>������<�2�!<"7�<�L��<`N<D��<��,�������N���?fff?��?&� ޔ@T�"!?��`?Uȩ?X�2!��z�!� Z��f/ǅ/�J�� �/�/�/�/?�/&??�J?\?G?�?��O%F ��o?�?k?�?W/O{)��?4O�8HmN H�[���G� F��=OvO�OsO�O�O �O�O�O�O___N_ ��o_yS;_���?�_O �_W_oo,o>o�So eo�_�o�o�o�o�o�oA��{�
r©{C�o ?�ocN}f��mtX����ç��}V{�BHP�\���Z܉r��p�q*�@I���}@n�@���@: @l��?٧]�� ��%�n��߱����=�=Dɋ�g����@�oA��&{C/� @��U���+J8���
H��>��=3H��_��� F�6�G���E�A5F�?ĮE��֏����fG��E���+E��E�X����>\��G�ZE�M�F�lD�
�� (��s�^��������� ߟʟ�� �9�$�]� H���l�������ۯƯ ���#��G�2�k�V� h�����ſ���Կ� ���C�.�g�Rϋ�v� �Ϛ��Ͼ���	���-� �Q�<�u�`߅߫ߖ� �ߺ�������;�&� 8�q�\������� �������7�"�[�F���j�����������(���4�����y���3�ϩ��<#q4 �{*<#q�0+#VhJ�jb��1E�䴛|���	�@� 6$�UP�	PhwQ�_���� ����� ���@1//A/g/R/#r$j/ |/�/�/�/�/�/�v_0??T?B<eZ?d?�?`�?�?�?�?�Q)�?��?OOBO0OfOtJ  2 H�6#v�H���C\�#vB�qqpB��p�pA#p@�O#t�s�O__�OC_�V�O�O�_��_�_�_�_#t^DR#p#p�!#p�F#u
 �_#o5oGo Yoko}o�o�o�o�o�o��o�o���Q ���R���4�$M�R_CABLE �2�R T�@�T~�A@� a?�ptq�Bmp��pʨ@B�@C�p�OM��`B�Xo�=�C�^��mjv³@·@B��@^M�O
�v�p��M7v�EC�kgЪ��x�@��@C��p9�t���uwZ*�v�[�����*�p�@��CL���r7�BV�9'�I`��sÏ �ޏ��ȏ-��6�(� "�P�F�X�������ڟ ��ğ)��2��q�Y&�������m�ү�����*�*�* FsOM ��Sy����]�7l%% 2345678901S��e� P���t�� �� j�A� �
z���not segnt ���WZ�TESTFE?CSALGRw0�D��Ad��Q��
(�u@�~�-rE��C�U�g�y� 9U�D1:\main�tenances�.xml����  � j�DEF�AULTK\FrGR�P 2�7�  �pRXk  �%�1st mech�anical c�heckz���Fd��l�u�vEE RZ�߲������ߜ<��controll�erL��e�:�wD���f�x�������MC���"8��� ����vEU�"�4�F�X�j���C������#���� $�6��CE�geA�.� battery:���vE	����������Sup�ply grea�sy1!B��8<B BIvE�v�К����N
caCbl5��
e :/L/^/p/�/I	�Y�/�)/�/?"?4?F?� $�/n?=�@��? �/�?�?�?�?
O Y?.O}?�?�?WO�O�O �O�O�OO�OCOUOgO <_N_`_r_�_�O;_�_ 	_�_-_oo&o8oJo �_no�o�_�o�_�o�o �o�o_o4�o�oj �o�����%� I[0�T�f�x��� ������!���E�� ,�>�P�b�����Տ� ��������(�w� L�������џ����ʯ ܯ�=��a�s���;� l�~��������ؿ'� 9�K� �2�D�V�hϷ� Ϟ��������
� �.�}�R�d߳ψ��� �߾�������C��g� y�N��r����� 	���-�?��c�8�J� \�n����������� )���"4F��j ����������� [0�f�� ����!�EW i/P/b/t/�/�/� �/////??(?:? L?�/?�?�/q?�/�? �?�? OOa?6OHO�? lO�?�O�O�O�O�O'O �OKO]O2_�OV_h_z_p�_�_\�B	 T�_ �_�_�__o0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p�����ަ�  �LQ?�w  @�A 
o ����F͏2�D�V���H*v�**  *Q(V!�������Ο��p���(���O_ HS��+�y�����_��� ӯ�/�A�S���?�Q� c���o��������� ���)�s���_�q� ��Ϳ߿������߀��%�7�Iߓϥ��J��$MR_HIST� 2�(U��� �
 \�B$ 23�45678901P�߼�~�p���9�O �%�����Om��� H�Z���������� 3�E���i� �����V� ��z���������A S
w.��d�����+��SK�CFMAP  �(U��"��� � 3CON?REL  ����\dEEXCFE�NB�
ZB�F�NC��JOGO/VLIM�d����EKEY��%_PAN�""�ERUN�+SFSPDTYP�<�DSIGN���T1MOT���E_CE_GRP7 1�(U\�� �P#��/��/"?�$? M??q?�?:?�?^?�? �?�?O�?�?7O�?[O mOTO�OHO�O�O�O�O �O�O!__E_�O:_{_�2_�_V[EQZ_E�DIT�$V#TC�OM_CFG 1��R��_o"o }
�Q_ARC_���%�T_MN_oMODE�&��Z�_SPLFo�UA�P_CPL�o�N�OCHECK ?�R *  �o�o $6HZ l~�������wNO_WAITc_L�'�W� NT�Q��RaU�<�_7ERR�!2�Rd� ��������j܏���a`Oj��q�|����_:��<9 � ?�?�Y�?��m,�c�PARAM:k��R�؆*��ܟǗf��� =  ��(�:�B��d�v�R� �����������ЫƗ��&�8�˟\�"ODRDSP�c�&��OFFSET_C�AR�PLo��DISܟ���S_Aa`AR�K�'�YOPEN_FILE���!%a�V�=`OPTION_�IO/!�M_P�RG %R%$�*O�a��WOް-��'كВ�\��  imr��M���	 ������	��r�R�G_DSBL  ���\U��o�R�IENTTO�f�C�l[A p��U�`IM_D��Yقr�Vv�LCT �F��R��%a��z�dj�_PEXi`�����RATig d��ԗ�UP )�{������(�X�L�Z��$��2�#��L�XL�pe���M��� ����������� �2� D�V�h�z��������� ������
�2��9 K]o����� �L�();M _q�����XY��.C�/+/X�P/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?2/D/�?�?�?�? �?�?OO)O;OMO_O qO�O�O�Ov?�?�O�O __%_7_I_[_m__ �_�_�_�_�_�_}��OƗ�*o<m��K��� ]ookQo�o�gmmK��o�o�g�g# +=[a��``����|҄�d	`���+���:�o�J�I�[�m��$�A�  ���o���؏ ��o���3��0�i��T���l�p�v�O��1������ ���r@ ����*�̐ @D��  ߑ?��ˑ?�5��5�D�  E�z����  ;��	l��	 ��@� �0��0� ��ې� � �� �U��H0#�H��G�9�G�ģG�	{Gkf�ˇ��o��,���C�?о�i��D	� D@ �D����r���  �5��>������B����� �BB�Bp{{�!5���O���bo�u�����Ӈ�����x�����(  ������׶���{�	'�� � �I�� �  �<��y�=���7�I�~��� <0��� � ?� ¯����������ҏ��z�NK���  '\���ġ� �C<�C�?�,�B���A������߰��@�����{�00ʉ��F�F���@5������� �������)��`�r�xT�d�5�� :�������x?�ff0�o���9� �p����� �85���>���ׇ��ʊΰ?�P�I�d�F�?�?���>�󙚋Ᏽ<2�!�<"7�<L���<`N<D��<��,w���������/�?ff�f?��?&���@�T�?�`�?Uȩ?X� )[�����ʉ�G �f��+����� ����+=( asJ���2T�V�/�HmN �H[�5�G� F��/W/i/T/�/ x/�/�/�/�/�/�/�/ /?яP?Z3?����? ��?8?�?�?OO�� 4OFO�?yOdO�O�O�O��O��\��B���KC�O _�OD_/]?���N_U_�_y_�çR����MD�HAХI��_�:hT�hPgQa�@I��@n��@��@:� @l��?٧�]�_ ��%��n�߱���=�=D�l��Hi��@�o�A�&{C/� �@�Ugo ��+J8��
H���>��=3H���_�o F��6�G��E��A5F�ĮE���o�`��fG���E��+E��EX��o��`>\�G�Z�E�M�F�lD�
��	�_T? xc������ ���>�)�b�M��� q���������ˏ�� (��L�7�I���m��� ��ʟ���ٟ��$�� H�3�l�W���{����� ���կ���2��V� A�f���w�����Կ�� ������R�=�v� aϚυϾϩ������� ��<�'�`�K߄�o��ߺ�ub(wa4����w����է�3��ϩ����na4 ��{��na�0+q#7�I�+�jbc��u�1E�䴛| ��������������x5P��PI�X1 e?r���~�����������������"H3nb$K]��� ����W?�5#e;E{i����)����#/�/G/U*  2 7H�6nfH���v#�\�nfB�A�A�@B)��P�PAn`@�O�/��/�/�/??(=~3 �R?d?v?�?�?�?nd��n`n`B1rn`c&ne
 �? OO(O:OLO^OpO�O �O�O�O�O�O�Omj�1� ��3����4��$PARAM_MENU ?����  �DEFPU�LSE�K	WAITTMOUTR[�RCVe_ �SHELL_WR�K.$CUR_S�TYLPP�\OsPT�!�_PTB�_��RC�_R_DECSN]P:�loo+o ToOoaoso�o�o�o�o��o�o�o,'QSS�REL_ID  ���W!�;uUSE�_PROG %�6Z%(�<sCCR�iPMrW!>S�w_HO�ST !6Z!�t��zTZ��s���q �:��{_TI�MEgRMv�u'PGDEBUGKp6[<s�GINP_FLM3SKc���TR����WPGA�� ��A?�ыCH����TYPE3\?0'!W� ��{�����ȟß՟� ���/�X�S�e�w� ������������� 0�+�=�O�x�s����������Ϳ߿ϔ�WO�RD ?	6[
 �	PR����MAI`��SU��QC�TE!����	9�TP�COL��lɴ���Lip ������ȵudw�TRA�CECTL 1�v��@Q G�_� 'G�U |����DT Q����$���D � �9�@U!9��0?��0?���?�P�0?��0?�=�=�=�=�=�1�CߨU�gߙ�	��
�����������C���C��C��C��C���C����Mp��*������u߇ߨ�߽߫�E��E��E*��E��E��E����w����}��� ��������������:� 
��.�L�^�p��#� 5�G�Y�k�}�������@��������Q cu������A cu������ �!�/�/�/�/�/�/`??1?C?U?-� u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� i?��ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/AS ew������ �+=Oas �������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_�oo)i�$PGT�RACELEN � (a  ���'`�=f_�UP ���e�lat`Xam`�=a_CFG ��leVc'am`���d�d�o�gO`�j�  ��e�bDEFSPD ��l�&aO`�=`H_�CONFIG ��leTc '`j'`d3t�Lb &a�6qP�d�aRq'`��=`IN�`TRL ���m�a8�egqP�Eu�"w��la�d2q�f=`LID�c��m	�yLLB� 1�"y 5�SuBBpB4��f Sx+�%�Vu�o << %a?�U�t�U�l����� ��ď�؏
�(�� �@B�p�V�x���Ú>� ڟџ��W�	�F�9��K�|��yGRP 1��|(a@� � �[�'aA?�x�D P�D�V�C2��$���7t�a���2q2p���p{�M��q�´L�.��BO�v�V�@��R���v���'a>'oY>a��ο���� =N�=R��W��Tύ�x� �Ϝ�6����ϼ�	�/��  DzT�]�'`
D߅�4ߕ߻ߦ��� �����'��K�6�H�@��l�������)(a�
V7.10b�eta1�d5p�B(�A�\)�A�G����>������Aw���*�ff��A�p�AgaG�����@�L���� ��o��������cAp��Ʋ�Bq�d ��#���²?���ߪffA����;�
oH3r&a �����6H2l�V�zKNOW_M�  �e�f�tSV7 �"zIrc� s�(:�^I[P�'a��sM���"{� ��	�e���x�t�d�������@�a�6!>%:/L,��V�qMR����T��h�Ƶ�/�+�OAD?BANFWD��s{ST��1 1�li�4pay�loa���>?)` �u)?n?M?_?�?�?�? �?�?�?O�?OO%O 7OIO[OmOO�O�O�O��O_�f72<�4>�O  �<I__���33_E_W_i_74 �_�_�_�_75�_�_�_o76,o>oPobo�77o�o�o�o78`�o�o�o7MA� ��0s�gOVL/D  ({���2PARNUM � ;�sS��SC-Hwy �u
��q8��#.�UPD��u�&�|�2_CMPa_�zp0� '�%~��ER_CHK�����!��������RS� �/��_MO��/�_��pe_REWS_G0�({
\� ���������՟ȟڟ ����/�"�S�F�w�j�]O�2PZ�j���O� �P��دݯQ��P��� �Q�+`7�V�[�Q�~` v�����Q��`��Կٿ�Q�$p����Q�V �1�5�!�@`�}x�THR_ICNR� |q��%d��oMASS�� Z���MN����MON_�QUEUE �P5�& ���pdN���UفN�����ENqD�9�5�EXEDߌ5�Z�BEC�%��O�PTIO"�B��P�ROGRAM %��%�R���?TASK_Iyt��OCFG ���x��� �DATA���)�@q� 2 @��L���������    �����"�t4�����  C��C�u��������IWNFO��m�� �����!3EW i{������ �/AS��������m�b�����K�_#��)����ECNBzp�sa�2���G#�2ʯ �X,		�=����6/��b%N!$�0�N)N)vě_E?DIT �)�/|�/�WERFLe��z��#RGADJ {̓*A�  5�? �5���&Ѫ���u�?�O  Bz�G �<N! ���%:r?�(�/#3f}2�/7��	HХl[�y�<1?O A�e��t$�6*z�0/�2 **:�2  ��?CM�u6B1E#���1;I�qa?]� [O)M�M9OKOyOoO�O �O�O�O�O�O�Og__ #_Q_G_Y_�_}_�_�_ �_�_?o�_�_)oo1o �oUogo�o�o�o�o �o�o	�-?m cu������ [���E�;�M�Ǐq� ��������3�ݏ�� �%���I�[������ ���ǟ�����w�!� 3�a�W�i�㯍���ͯ ïկO����9�/�A����e�w�������r�	 <�F�� 4�m�X��9�π�3[ϼ�W�����7P?REF �/:~��
�%IORITY��ך&��!MPDSaP���*W2M�UT�|�3�&ODUCT���*�ϛ6OG�0_TG� �*���HIBIT_DO��(��TOENT �1ѓ+ (!?AF_INEw�*�~5�!tcp5�>]�!udL��?!icmt�{>֌�XY(3ғ,��!)� 	A����� ���$���P�7� t�[�m�����������@��(L^*��(3�/9W2`?���3�>b���	G/�L��4��8�>A~Q2,  �%Ѐ�N`r��%�6�Z������3�sENHANCOE ��2A�Ad�Z/A%������(��!�!PORT�_NUMx�� �D��!_CART�REPX����SK�STAw���SLGmS'�����Q3�^�Unothingb/??Q?c?��0TEMP ؛��o?�'0_a_seiban���?�� �?O�?,OOPO;OtO _O�O�O�O�O�O�O�O __:_%_J_p_[_�_ _�_�_�_�_ o�_�_ 6o!oZoEo~oio�o�o �o�o�o�o�o D /hSe���{9�VERSIVЙ���p disa�blet"w;SAV�E ٛ�	2670H755�x	�O�!J/Q�c��� 	�����݋ԏ�e��,�>�P��^�	�������_��� 1���<��Ԑ �ѵޟ�ͷ�URGE B���޿�WF���z�4"��W�#�=�bѹ*WRUP�_DELAY ���-��WR_HOT %+Ƅ�I/���N�R_NORMA�L���Ҭ��ЧSE�MI��E��QS�KIP��܆'͓x ��������ҿ��#� �1��+�=�O��s� aϗϩϻρϓ����� �'�9���]�K�mߓ� �߷�}��������#� ����Y�G�}���g�����������R�BTIF>���9�C_VTMOU�'�%��9�DCR��޾h� С�B��4Bu >�-�G:Q%��jp����J���������<2��!<"7�<L���<`N<D��<��C����I[J���� ���!3Ey7�RDIO_TYP�E  Ý;QE�D T_CFG ��$-U�BH%�E��b�2�$+ �8BȖ��*8 */��N/9/r/]-/�/ 2��/��/���/�/? E?3?i?W?�?w7�/�? C��?�?�?O�?/OO ?OAOSO�O�?�O�?�O kO�O_�O+__O_=_ s_�O�_�Ok_�_g_�_ �_oo%oKo9ooo�_ �o�_woQo�o�o�o �o5#Y{o��Q �M�����1� �U�w|��]����� ӏ������	�+�a����x�E�INT �2៩����G;� ��ț"5�b(f�0 � �=�@� 1�P�R�d��������� ί�����<�"�4� r�`�������̿��� ޿��8�J�0�n�\� �π϶��Ϯ������ �� �F�,�j�Xߎ�+��EFPOS1 1��n  x f��ٻ����)�5� �����|�g��;��� _���������B��� f������7�I����� ����,��P��M �!�E�i� ���L7p� /�S���/� 6/�Z/l///S/�/ �/�/s/�/�/ ?�/? V?�/z??�?9?�?�? o?�?�?OO@O�?dO �?�O#O�O�OYO�O}O _�O*_<_�O�O#_�_ o_�_C_�_g_�_�_�_ &o�_Jo�_no	o�o�o ?oQo�o�o�o�o4 �oX�oU�)�M �q�����T� ?�x����7���[��� �������>�ُb�t� �!�[�������{�� ��(�ß%�^������ ��A�ʯܯw���ï$� �H��l����+���xƿ_���2 1�� h�z���2��V�\�z� Ϟ�9ϛ���o��ϓ� ߷�@�������9ߚ� �߾�Y���}���� <���`��߄���C� U�g�����&���J� ��n�	�k���?���c� ����������	j U�)�M�q� �0�T�x %7q����/ �>/�;/t//�/3/ �/W/�/{/�/�/�/:? %?^?�/�??�?A?�? �?w? O�?$O�?HO�? �?OAO�O�O�OaO�O �O_�O_D_�Oh__ �_'_�_K_]_o_�_
o �_.o�_Ro�_vooso �oGo�oko�o�o�o �o�or]�1� U�y���8�� \�����-�?�y�ڏ ŏ����"���F��C� |����;�ğ_��ο�3 1�뿕��� �_�J�������B�˯ f�ȯ���%���I�� m���,�f�ǿ��� ��Ϫ�3�ο0�i�� ��(ϱ�L���pςϔ� ��/��S���w�ߛ� 6ߘ���l��ߐ��� =�������6���� V���z���� �9��� ]�������@�R�d� ������#��G��k h�<�`�� ���gR� &�J�n�	/� -/�Q/�u//"/4/ n/�/�/�/�/?�/;? �/8?q??�?0?�?T? �?x?�?�?�?7O"O[O �?OO�O>O�O�OtO �O�O!_�OE_�O�O_ >_�_�_�_^_�_�_o �_oAo�_eo o�o$o �oHoZolo�o�o+ �oO�osp�D��h������4 1������� w����ԏo������� .�ɏR��v����5� G�Y�����ߟ���<� ן`���]���1���U� ޯy����������\� G������?�ȿc�ſ ����"Ͻ�F��j�� �)�c��ϯ��σ�� ��0���-�f�ߊ�%� ��I���m�ߑ���,� �P���t���3�� ��i�������:��� ����3������S��� w� ����6��Z�� ~�=Oa�� � �D�he �9�]��
/� ��/d/O/�/#/�/ G/�/k/�/?�/*?�/ N?�/r???1?k?�? �?�?�?O�?8O�?5O nO	O�O-O�OQO�OuO �O�O�O4__X_�O|_ _�_;_�_�_q_�_�_�o�_Bo(�:�5 1�E��_o;o�o�o�o �_�o%�o"[�o �>�bt� �!��E��i���� (���Ï^�珂���� /�ʏ܏�(���t��� H�џl������+�Ɵ O��s����2�D�V� ���ܯ���9�ԯ]� ��Z���.���R�ۿv� ����������Y�D�}� ϡ�<���`����ϖ� ߺ�C���g���&� `��߬��߀�	��-� ��*�c��߇�"��F� ��j�|����)��M� ��q����0�����f� ������7������ 0�|�P�t� ��3�W�{ �:L^���/ �A/�e/ /b/�/6/ �/Z/�/~/?�/�/�/  ?a?L?�? ?�?D?�? h?�?O�?'O�?KO�?xoOUogd6 1�ro O.OhO�O�O
_O._ �OR_�OO_�_#_�_G_ �_k_�_�_�_�_�_No 9oroo�o1o�oUo�o �o�o�o8�o\�o 	U���u� �"���X��|�� ��;�ď_�q������ 	�B�ݏf����%��� ��[������,�ǟ ٟ�%���q���E�ί i�򯍯�(�ïL�� p����/�A�S���� ٿϭ�6�ѿZ���W� ��+ϴ�O���s��ϗ� �ϻ���V�A�z�ߞ� 9���]߿��ߓ��� @���d����#�]�� ����}����*���'� `�������C���g� y�����&J��n 	�-��c�� �4���-� y�M�q��� 0/�T/�x//�/�O�D7 1�OI/[/ �/?�/7?=/[?�/? ?|?�?P?�?t?�?�? !O�?�?�?O{OfO�O :O�O^O�O�O�O_�O A_�Oe_ _�_$_6_H_ �_�_�_o�_+o�_Oo �_Lo�o o�oDo�oho �o�o�o�o�oK6o 
�.�R��� ��5��Y���� R�����׏r������ ���U���y����8� ��\�n�������?� ڟc�����"�����X� �|����)�į֯� "���n���B�˿f�� ���%���I��m�� ��,�>�Pϊ������ ��3���W���Tߍ�(� ��L���p��ߔߦ߸� ��S�>�w���6�� Z��������=��� a���� �Z������� z���'��$]�����@��/�$8 1��/v��@ +dj�#�G� �}/�*/�N/� �/G/�/�/�/g/�/ �/?�/?J?�/n?	? �?-?�?Q?c?u?�?O �?4O�?XO�?|OOyO �OMO�OqO�O�O_�O �O�O_x_c_�_7_�_ [_�__�_o�_>o�_ bo�_�o!o3oEoo�o �o�o(�oL�oI ��A�e�� ���H�3�l���� +���O���ꏅ���� 2�͏V����O��� ��ԟo��������� R��v����5���Y� k�}�����<�ׯ`� ���������U�޿y� ϝ�&���ӿ�π� kϤ�?���c��χ��� "߽�F���j�ߎ�)� ;�M߇�������0� ��T���Q��%��I����m�����MAS�K 1�����:�H��XNO  �)�G�M�MOTE�  i�  ��_?CFG ������PL_RAN�G�������OW_ER �� �SM_DRYP�RG %�	�%���S!TART ��a
UME_�PRO0B��_�EXEC_ENB�  ����GScPD� � ��gTDB�RM�IA_OPTI3ON���� ��INGVERS`�j���I_�AIRPUR�� ��
w���MT_�"�T ��OBOT_ISOLCg��������%NA�ME����OB�_ORD_NUM� ?��H755  ���/�/�)�PC_TIMEOUT��{ x�S232���1�j� L�TEACH PENDAN� ����64h,����Maintena�nce Cons���3?U6"O?��?No UseC=? E?�?�?�?�?�?��"GNPOp �"��n��!CH_L� �� .��	nA9O!�UD1:�O;OR�!�VAIL�!d������SR  ��l��GER_�INTVALc���P]�IV_D�ATA_GRP �2�j���� DPP��_��_�Y j��_�W�_o�_+oo Oo=o_oaoso�o�o�o �o�o�o%K9 o]������ ���5�#�Y�G�}� k�������׏ŏ��� ��/�1�C�y�g��� �������ӟ���	� ?�-�c�Q���u����� ���ϯ��)��M��;�]���q���n��$�SAF_DO_PULS��o�8A��ѱN��CAN�"c���A SC ���`XW����
>!����!~1~5!���  �_Y�k�}Ϗϡϳ�Bπ��������1�,H8C��2Z�!�eّdZ�uі�	�<� @���߻����։��� P���_ @��Tl��4��F�X�e�T D��e���������� ����0�B�T�f�x��������OE���������  =/5;�o_4-�Qp*U/E
�t��Di� ��1�
?  � �0*1� )�������� ,>Pbt� ������// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6?H?Z?l?�1��ߕ?�? �?�?�?�?OO%Ot? H�QOcOuO�O�O�O�O@�O�O�O�A5O��0�� M�D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����?8�J�\� n���������ȏڏEO ���"�4�F�X�j�|� ���O'U1_��Ο��� ��(�:�L�^�p��� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/πA�S�e�wωϛ�p� ��t��������+� =�O�a�s߅ߗߩ߻� �����������\G�Q����@��	12345�678fh!B�!��������,����������� �#�5�G�M���p��� ������������  $6HZl~�� _�����0 BTfx���� ����/,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?�^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O O?�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�O
oo.o@o Rodovo�o�o�o�o�o �o�o*<�_` r������� ��&�8�J�\�n��� ��Q��ȏڏ���� "�4�F�X�j�|����� ��ğ֟�7���
�����A�S�e����Cz  Bp�� �  �r�2��� } �r�
���  	Ĥ������ �/�	��0��دu����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��Z�����%�7�I� [�m�ߑߣߵ����� �����!�3�E�W��<�0�̡p�<�����y�̡  �����_��ССt  ������_��`<��$SCR_�GRP 1��*P3� �� �<� �k�	 7��?�P�I�1� q�`�_�\���x���u�g�����C������E�V�����S��LR Mate� 200iD 5�67890ΠL�RM- 	LR�2D 4 9�
1'2343��>�7��� �?���.� ��.�S����M����		���%~5��H�?��C�.�fu�v��}���<����p/h�+�� h��_,X�_JE�[�Bǈ��a/_"x$[�9A���/  @<��%f[�@�� �/ ?����%["H���/�*[�F?@ F�`2
? /.??R?=?b?�?s? �?�?�?{�_!�!�"�?0�?�?
ODB�*O�? pO[O�OO�O�O�O�O �O_�O6_!_Z_D�jZ ����W�_k����_��_<��!@��>�A�j�_}�@� o���5gYY���uo�9�A� �V�e��$�`S�u<� �o�o�oz�ax#5	.�\s
��i{��T_���9��EC�LVL  <������`Q@�qL�_DEFAULT��tJ����<��HOTST�R��a�qMIP_OWERF�p}��#�L�WFDO�� #��rRVENT� 1��q�qD� �L!DUM_E�IP����j!?AF_INE�܏�9�!FT����ҏ/�!bT� ���{�!RPC_OMAIN|�^��j��ǟ��VIS���������!TP�P�U
�ŉd�_�!
�PMON_PROXY`�ȆeN���&��y���f����!R?DM_SRV��ŉ9g�C�!Ra_��ƈh2���!
��M�¯i~�ۿ!R�LSYNCܿ��8ʿ'�!ROS̱�N��4�s�!
�CE(�MTCOMdt�ȆkbϿ�!	��OCONS��Ǉl����!��WASR�C�Ȇm��W�!N��USBX�ƈnF�>��!STMx���Ċo����B��������<�a�(�� ���*SYSTEM*�wPV9.3044� ��1/9/2020 A �zPܝ��� y���_S�PD_T[����_TRQ  � 
��AXIS��� ���� �2x ��DETA�IL_  l�$DATET�IME{P$ER�R��DC�IMP_�VEL   �	U�TOQ]�AN�GLES]�DISyTg���G_NAB��%$L{�D������REC�� ,� ���!�2 $M�RA�� 2 d��IDXD����� c`$OV�ER_LIMIT�]� 	��OCC�UR��  �H�COUNTER���FZN_CFG��� 4 $EoNABLC�ST=��D�FLAGD�DE�BUaRv� �4GRf�  �� 
$MIN_�OVRD{P$I�NT_r���F�ACE�SAF>�MIXED��	��ROB��$�NE�PP��HE�LL; w5$J� BASC��RSR_I  �$N��1]� �01��12T3�T4T5T6T7rT8��$ROO�������T_ONLY�{P$USE_A�BO7��1ACKgENB\��IN���T_CHK�OPq_�T �_PU��'M_@�O.�E�PNS4���T ��MN�TPFWD_�KAR[��I�RE=P�OPTI��E�QUE;)��DV"Y�
$CSTOPIg_AL�EX���� C�XT M1b�)2D�� TY��SO� NB�DI��TRIa�!['I�NI����#NRQ�06� END4$�KEYSWITCaHB#W!1�$HEX �BEATM�#PE�RM_LEZ�b!E�W��7UV#F�$W"SV4DO1�M� O
�EFPS����b�5� %C�0��E��OV_MS!R E?T_IOCM���2d�&�!xHK�	 D H�1S�UB�"MP�I�P�O�$FORC�A#WARN#LOM�*  
 @;@F�U���SU��5!A�R� �E2�F3�F4��A���Og L�B<��<(UNLO @���DED@�(��S�NPX_AS>; 0?ADDq s�$SIZC�$�VAR��M�IP��S�@A�A � $,)P�2C	APD�BCV�VFRIFD���SЇ �I�4)�F34OD?BUS_AD/A��S�Y{$' ML1DI�AxA$��MY1��!e3h4a�S|2 � 0P�s�TE
d8bS�GL>aTA@  &S WcB��P`�?`��T�!pcPSE�G�"paBW� @dS�HOWxeE�BAN��`TPOF�Qd9�h0h�!��VCڜ G� L`$P�C�����`��$FBX�A���fSP� A���e�aD�`�7� �;�A0��K }�?q�@Fw�@Fw�@FwT�@Fw5Dy6Dy7DyU8Dy9DyADyBDy@�@Fw �Fw�`FwFDx �`�Py`�jy$`���y1�y1�y1�y1��y1�y1�y1�y1
�y1�y1���هPyU2]y2jy2wy2�yU2�y2�y2�y2�yU2�y2�y2�y2�yU2�y2�3Cy3PyU3]y3jy3wy3�yU3�y3�y3�y3�yU3�y3�y3�y3�yU3�y3�4Cy4PyU4]y4jy4wy4�yU4�y4�y4�y4�yU4�y4�y4�y4�yU4�y4�5Cy5PyU5]y5jy5wy5�yU5�y5�y5�y5�yU5�y5�y5�y5�yU5�y5�6Cy6PyU6]y6jy6wy6�yU6�y6�y6�y6�yU6�y6�y6�y6�yU6�y6�7Cy7PyU7]y7jy7wy7�yU7�y7�y7�y7�yU7�y7�y7�y7�yE7�y7����`P�0=U�� �����I
���R x? $TOR�!�P  _�MO����6��Q_ RE"rn�(�b@]�S�CX!(�B�_U�PM�xY�SL�� � 0U�RN�T%We ?px�0y�
rVALUN�	 \&��Fj�ID�_L33��HI��I~xB$FILE_0#����$�3�@h�S=A�� h��1�?E_BLCK�#>�|YaG�D_CPUW��1PW�%PY��PY�d`*#R  � PW ��P��LA~aS��������RUN_FLG ��������Z0������H* ��' ��PQ�T2\!_LI�B�  #G_O��"d P_EDI��(`T2� G�O�I�R�xP�P ��TBC20t ��5`���P�GFqT�$��#TDC��A1^ � M�P��&�TH�PnQ���R� PI@ERVAE�#*�#*a����  X ;-$ULEN�#b�#U� RA� �Bi��W_#��1U��2&�MOO��ES�P�I >������U��DE��QLACE�B�CC�C>�0_�MAP�"%�"!T#CV),J!�T<1K* j%`*r�q�%�q�J� AuM�$�0JH"7.p��!�a�2�0�P&p�!� PJK 6VK�a1a1�a0J�a*13JJv3JJ&3AAL3@L03L0F6%aJ25} N1q,}0<+& <�L�_la�0�ќ C�FR `��GRCOU��Za�RqN� �CnS�0REQUI9R�PEBU�SQn�&$T�2A�R�6�P� \��@�APPR@C�L<�
$X NKHCLO� [IS�pI��
�YV � M�� ' | �B�D_MGa�@C0p2�Hp$ ��GBRK�INOLyD�F�`RTMOFHZ�M�EJF  TPN4  3 &3 j3 s3J 6;U7;ULac�|Q�� B�|�a�Wa�SPATH�W�Q�S�Q��S�@@@��`SCA��WLB�AINTU�C��`CpUMhY���� $a���0?j�P?jK?`PA�YLOA�GJ2L���R_AN��cL����i�azi�a�ER_?F2LSHR$�aLO�dba�g!c�g!cACRL_�ep�grdt2H��<�$yH�B2rFLEXNCu�J� P8B@��);�0OJT :as� �w�tvu1���F1�q)�=������/m�E/(/:/ L/^/p/�/�/�/D�a� �'�# 4Q�s��/�/�/$�q�*T��B�X*�K� �%����	5��?'? 9?K0O5X5F5j5s?�?ؗ?�:m BJ�4  ��� �?�?�?�0��A1TV� A� ELĀ�(�HJ@@JE��@CTRaQ�TN���$��7HAND_�VB<�Nq���T!� $��F2�F�ƭ�SW�1�S�F"� $$M�`�I� �Aո�A��ص)RƁA��w`�F�� ɸMA(�L���JA�KA�K+���Kp��JD�KD�KP2�PG����ST�G��4�I��N�HDY��I@ �F�3Ř`V�g�q�g��ayg 7�����EP CULUUU^UgUpUyU�R:�2J�# ˰�t��R ~���}A��A'SYM�U>�@�V!"/�l�ao_& �h `,d]䜸6oHoZolo~cJ�l6P�j���\�ic�_VI���<}C�V_UNf���;��aJ52�`�2� �l6��eC�g��m� y 6P)���?tGs�M� HR� �$0����ap[DI�@�3�O�2��ӣ% K�:�I�A:Q�c4 W�B�BZ�4��Pǀ�� & � ��ME����]��D�T��PT�๠�P��0Ť`p|����	�T��1 $D�UMMY1K$7PS_T�RF��0�$��@FLAƾ0YP���$GLB_Tΰ���� iq�0��U�a' �X8@�7�QST���@SBR�PM21�_V�"T$SV_�ER�`Oo�[sC)L/[AŀO7���GL��EW�1( �4�0�$Y��ZB��W�� �a��A^ �b���U�) �N���$GI�e�}$� �(Π���1* L��0�n�}$Fn�E^&NEAR��N[�yFH)��TANC[�����JOG
��,P +ˠ$JOINT�������MSET�1,  "�E.%Ɓ�S���P�"�1-�  �]�U��?�@LOCK_FO�`�� oBGLVX�GL�(TEST_XMN@N�!EMP� k�2-� $U�p���#2)@�<1*2��4� <1(]CE�0
#�]0 $KAR�M>	TPDRA�z4�q!VEC�p�6u I�U<1+A1HE� T�OOL��3V�R�E�0IS3�u�26�^QQ�ACH� @,��1O�P��3�Q�	 SI>B  @�$RAIL_BO�XE���ROB�O4?��HOW�WAR:q,A� �1ROLM�RE���4cBp�@E��PO_F��!�HTML5��a������Ҡt�1�Q.}/ �R�0�O�r/�B��!�@v�OU�"0 t��85(D�.��� RPuO�A�PIP6N���2B�1c�<1�@~�pCORDED� ��P�@E XT+P�)�P�OD  1o D OB`� 2�� �WzQ�zRn��4�SYSzQADR�3���� TCH� o2 ,��EN��*jqA�!_��T�����VWVA`3 � �0���PREV_RTmѿ$EDIT,fV/SHWR�GK`������Do 3��bd;�$HEAD���|`��4cKE|�� CPSPD�f�JMP�PL��
�3TR��4�P_q��VI0S3�Cy�N�E�04�o�TICK����Mhq�ҽcHN=5 @�P�ať��a_GP*vFkpS3TY�R�1LO/�P�p�b&r�p6�@
'`MG�U%$a�=GS)�!$(���t� 1 �P
�*vSQ�Ut0���TER�C� ���SӤ7   S槤��t�ħ1�O� }_�IZh���PR]P0�H��a�@PU��X�g_DOM"�PXS� �K��AXIw�vCA1UR�Ń4�3@pȥV���_�0�RET���P�"�P��vpFd��wpA������9 G2K�"SR��8l�pι� ݺ3��E��3��3� �3�,�y�N�y�^�y� nƋ����ɋ�ɜ�ҩ�	C���Cȝg�y��ܝ��SSC 79 h�DS8p{1f� SP. ��AT\���Y�p�b�AD�DRES�3B7`S�HIF�B21_2C�H3��QI6����TU6I� :>�BCUSTOل��V�"I";�R�(��T<���
:
��V�A�h�b < \EX� vpG�� `��C����܂V�Vy���TX_SCREE|R=��=�qTINA� �״��Q������> T�av<��QuR�$ƅ��R�� �3`RRO7�b �P�`�Sa;UE�d? ����Qr� S��QRSMp�{�UfP�p������S_���!������!�⹁C�"��� 2->ҰUE��@(�\��H�GMTz�LT����b"Q�"�B�BL_�0W� b AS �vpN�O�Z҃LE�e�2@�d�RwIGHn�BRD��ߡCKGR� ��T�gP�ג�WIDTH� CX`R���17�UI�@EY�@aB d��@Q@Zr@=D�BACKXq�4	�h FOTQ�LABc�?(h I<�0�"$UR8AI�� ��n HD� C 8��b _{a��l�o R��"� H�n RY�O�b D!p����Uzк�R�"]AL�UM�㜆٠ERVHQd���PL ��Ef �GEM�3!׀mR&�`LP��E�pj�))�z�7���7��06�U54�64�74�8��r%�C�L ����1��!S `D��US=R�F <En 1U�,��FO��PRI��m@&� �TRIPAm�oUNDO�dG���p$ }�DA|���832���p Hg���.G�G �pTv@X�L��bOS�wR��J�N�1>I�����:t�32U�>J������9uNOF�F0�K���O- 1I P?-J PGU�QP>�"pZU�d��SUB:r� vrE_EXE��PV�aNWON� �L� n��WA�7`��1�ՠV�_DB���Q��T�� �M!ra!�@'�O9R�0 %RAU,�$�T)�W�_*`�dNs |5��XOWNQ >�T$SRCU����pD0l%*�MPFqIQt����ESPT� ���5��A���2M8<"E`�O `� �r�T��pCOP�$��S _� �2�!�A5�CT�Ӧ�#���2�`PB/� �P�SHADOW����3P1_UNSC�A�3P3��]3DGD<�1�QEGAC�#<���QPG۲Q (��NO���LpPE�����VW�4cqG|Ā�R � �P�VEU���2ANG����6�6��2LIM_X�%F�%FH *AL���7 ��0��VF��#�VCC�zp�dS�2C�pRA�|w�0�u�bNFA�2`5pE�Q2 G����RRS �DE�2���STE a�3��ܣ�!��Y4� �;�)A�s� �1+U�PP_AFP�C�@[��@�T� Ar�Q�sA�El]�q��/�C���mUDRI�0lV�1V�3p�T�`+�D��MY_UBY���M��uV��p�ia�X41
b�P_f0�$bL^�B�Ma�$�`DEY��cEX'Qu6QMUj�`XWM��US���� _R�����z�6G�PACI�D �0v!�4�b�b��b���RE���g8RS�bpU �� �G�0P���`�SSR� ppV�г�C��ъi	�"u�RTSW�` �Ci�0caF�O����A�hs3�E%�UEd�3id�SSHKZRW���z�1+�ep)��3EAN�y��hu�� SRMRCV�X� ��O�@M�C»�	�r�c�rREF:����qB�?p ���zP��P��r���_i �z���{�� P a�C��R˰�B�SR�Y ��1��5rܣ��~�U$GROU�� ��c(��C�@T
uY��2��$ذ��e 0��V��Y�<��٠UL��AW� C6@��XR`O�NT�#��42�� �᜖��[�Lcŕ@cŕ��ї��AT!�nq�Z t� MD��HPHU�A�0�SA.�3CMPU�F�0�(��_��R�D��P��sЁXc��1VGF|?0r�[, &��qM���PUF_S�01b�`0�ROx�,��;��U��L�SbUR1E����bRI�c�IN�#��?
OKt!�.It!�qGINUbH��H��V�=B�Q���ӥ�WW�gQ�S6Sa�yfLO@�S�1pP��U���NSI�D��!0�4��4�>HX�_PE=�Yg�Z_IM-S�2W�Ys4C�2���R�ǂ�RSLN/\ �"�?1M R���UaCG`GtA �P�l�r�v� ��!e ��h����į֯�N���o��~� �`IA�] ��HDR���JO��"��$Z_UP+Q=�_LOW�վ�tZ�t��2LIN�EPO��o	�Ѿ������A�D��gR���^ 5h�PA�THc  h�CACH��m�
�����u1T0�#C9AIT�F���TD���$HO��Rr����S��v���������!PAGE�� VP�b�@8�O_SIZ�CB�ZCP`=�+S@���CMPb���AIMG�4	�A9D���"MRE���G�GPPH`� 6A�SYNBUF6V�RTD����G��DLE_2D=Dɲ	%C�AUAc
�Q�p���ECCU�hVEM��`m�T��VIRC����������LA|�c�!NFOUNo��DIAG 	RUaX#YZ��UaW%q��H���q T�@BbI�M��u0��GR�ABBցYSqpLKERz`CD�߂FS�=��50D͑GۑS4R���_�pppCKLAS��|qR���`  W��T$�c @�R�T$R��@��a �1�� u���Ti�!XQ� ���e�I�J���B9PE3VE�A�PPK�`�l���GI�NO�!�Ba�q3pHO� �Bb � b���H�� y&S���7�"RO>�3ACCELO�MQ-�%VRo�UG�� ��!Bb�0& AR�3P�A� �.[�D�3RE7M_B� �@3p�JMh�&rc���$SSC��{�3p
����0d ��
�S���Nc4�pLEX��e T�ENA�B�Bbg�CFLDR�HFI �G���H�8d�s� C�VP2>X�f� $���V�a�MV_PI �C�4H�P�@�P%�I	F�/RZJ;D3E@`H�$HH�3E�1GAREΥ�LOOS��JCqB�J'2�CON8�SPLAN� ��"�C�F+Ut/�)I��GM pa�KTUFS�PUa �E+QH��EgG�-�4 dLRH��!< RKx�!VANC�3��Rs_O���0g (��=�L��c#$Һ�Rs_A?@�0h 4���_�^p� n�O�&ri� h~p+9��n��OFF, ��g� �� ���EA%�
��< SuK��M`�VIE�`2h �P��0�j < �:脯Ԣ������pD�@}���CUST���Upk $W�T�IT-�$PR�l1�OPTqlq��VSF�p�l�� �p�	��1SMEO��mY2�3�$J�`�؅�u�_g��`n�Y2�g���_���X�VR��o}�`T��%�ZABC��p �r胺9�
���ZD4 CwSCH�q L�` �t� �
�5�!��ӀG�GN)��rLu���p�_FUNX��� ���ZIP��r,Y2# LV<�L₎���`�ZMPCF��usrU��r�!h�D�MY_LNX`Ma �T����tt �$����m�CMCM���C<�C6���-�P~�Q $Jǃ��D-�͂ނׇېㅄې��_��<�܂�U�X�l�UXEUL -��҅&��&�8�J�x8�Z�ƀFTFLʆ܇�/��Z+�u� :{F���p+�Y��D v 8/ $R��U�AN��EIGH�#�h?(�(0yv�qœuw a�q �c,��p$B����Psb_SHIYFT�=xRVf Fsp&�p	$E�� C��@6�d�`Ұ�1r�
�4���D��TR��puV�QC��SPH� ��x ,(0ܘ����$G�I��KL ?%�����  �(%SVCPRCG1�`*�5��25�D:�$�3]�b�$�4��D��$�5����$�6տDڿ$�7���$�8%Ϥ*�$�9M�R�!�0 u�{�%�'���$�O��� $�w���$����$�ǿ B�$��j�$�ϒ�$� ?Ϻ�$�g���L���
� L���2�L���Z�L�� ��L�0ߪ�L�X���L� ����L���"�L���J� L���r�t� ����$� ����D�* N9r]���� ����8#\ Gn�}���� ��"/4//X/C/|/ g/�/�/�/�/�/�/�/ ?	?B?-?f?Q?�?�? �?�?�?�?�?O�?,O�O>ObOMO�O��݀V� ���M{C:�H4���D�� 2���`��bx 	���,���O	_R�O2__ V_=_O_�_s_�_�_�_ �_�_
o�_.o@o'odo Ko�o�o�O�ouo�o�o �o�o<N5rY �}������ &��J��o?���7��� ��ȏڏ�����"�4� �X�?�|���u����� ֟��ϟ�c�0�B�)� f�M���q�������� ˯���>�%�b�t� [������ο%�򿩿 �(��L�3�pς�i� �ύ��ϱ��� ���$� �H�Z�A�~�տsߴ� k��߿������2�� V�h�O��s����� ����
����@���d� v�]������������� ����<N5rY ������Y� &�J\C�g� �������4/ /X/?/|/�/u/�/	 �/�/�/?�/0?B?)? f?M?�?�?�?�?�?�? �?�?OO>O%O7OtO.{Cd �{F	bO�O��O�O�O�O�O_&[%��&_K_RS��� dQQdUt_�Wl_�_�_ �_�_�_�Y8_o`Y�_ Jo8ono\o~o�o�o�o 
o�o.o�o"F4 jXz�o�o�� ����B�0�f�� ���V���R�Џ��� ��>���e���.��� ������̟����X� =�|��p�^������� ��ȯ�0��T�ޯH� 6�l�Z���~�����ۿ ��ƿ���D�2�h� Vό�ο���|����� ����
�@�.�dߦϋ� ��T߾߬��������� �<�~�c��,��� ���������D�j�;� z��n�\��������� ���@���4��D jX�|���� ��0@fT ����z��/ �,//</b/��/� R/�/�/�/�/?�/(? j/O?a??:??�?�? �?�?�? OB?'Of?�? ZOHOjOlO~O�O�O�O O�O>O�O2_ _V_D_ f_h_z_�_�O�__�_ 
o�_.ooRo@obo�_ �_�o�_�o�o�o�o *N�ou�o>� :�����&�h M�����n������� ڏȏ��@�%�d��X� F�|�j�������֟� ��<�Ɵ0��T�B�x� f���ޟïկ������ ��,��P�>�t����� گd�ο��޿��(� �Lώ�sϲ�<Ϧϔ� �ϸ�������$�f�K� ���~�lߢߐ��ߴ� ��,�R�#�b���V�D� z�h��������(� �����,�R�@�v�d� ������ ������� (N<r����� b����$ J�q�:��� ���/R7/I/ / "/�j/�/�/�/�/�/ */?N/�/B?0?R?T? f?�?�?�??�?&?�? OO>O,ONOPObO�O �?�O�?�O�O�O__ :_(_J_�O�O�_�Op_ �_�_�_�_o o6ox_ ]o�_&o�o"o�o�o�o �o�oPo5to�oh V�z����( �L�@�.�d�R��� v����� ��$���� �<�*�`�N���Ə�� ��t���p�ޟ��8� &�\�����L����� Ưȯگ���4�v�[� ��$���|�����¿Ŀ ֿ�N�3�r���f�T� ��xϮϜϾ��:�� J���>�,�b�P߆�t� ������ߚ���� :�(�^�L���ߩ��� r����� ����6�$� Z������J������� ������2t�Y�� "�z����� :1�
�R� v����6� *//:/</N/�/r/�/ ��//�/?�/&?? 6?8?J?�?�/�?�/p? �?�?�?�?"OO2O�? �?O�?XO�O�O�O�O �O�O_`OE_�O_x_ 
_�_�_�_�_�_�_8_ o\_�_Po>otobo�o �o�o�oo�o4o�o( L:p^���o �� ��$��H� 6�l������\�~�X� Ə��� ��D���k� ��4����������� ��^�C����v�d� ������������6�� Z��N�<�r�`����� ����"��2�̿&�� J�8�n�\ϒ�Կ���� ����~���"��F�4� j߬ϑ���Z��߲��� ������B��i�� 2������������ �\�A���
�t�b��� ��������"��� ����:p^��� ���� "$ 6lZ����� ��/�/ /2/h/ ��/�X/�/�/�/�/ 
?�/?p/�/g?�/@? �?�?�?�?�?�?OH? -Ol?�?`O�?pO�O�O �O�O�O O_DO�O8_ &_\_J_l_�_�_�_�O �__�_o�_4o"oXo Foho�o�_�o�_~o�o �o�o0T�o{ �Df@���� �,�nS�����t� ��������Ώ�F�+� j��^�L���p����� ��ܟ��B�̟6�$� Z�H�~�l����
�ۯ ������2� �V�D� z������j�Կf�� 
���.��Rϔ�yϸ� BϬϚ��Ͼ������ *�l�Qߐ�߄�rߨ� ���ߺ����D�)�h� ��\�J��n����� 
���������"�X� F�|�j���������� ����
TBx �����h���� P�w�@ ������/X ~O/�(/�/p/�/�/ �/�/�/0/?T/�/H? �/X?~?l?�?�?�?? �?,?�? OODO2OTO zOhO�O�?�OO�O�O �O_
_@_._P_v_�O �_�Of_�_�_�_�_o o<o~_couo,oNo(o �o�o�o�o�oVo;�zo�a�$SERV�_MAIL  �ezp�`xOUT�PUTox��`@dtRV 28v�`}p (qJ<�dtSAVE�|~y�TOP10 2>�y d �o6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я����0�*�u�YP�as�FZN_CFG ;u}s�t��q�uj�GRP 2�t�� ,B �  A���aD;�� B���  B�4�sRB21��vHELLm�u�v�p����,�%RSR,�-�?� x�cϜχ��ϫ����� ����>�)�b�M߆���ߪ��  ��zҪ����߸��� b�`�������
��2�`d��U�߶�HK 1	� ��������� ���.�)�;�M�v�q��������������ټOMM 
�-޲�FTOV_ENB�ot�q�um�OW_R�EG_UIMbrIMIOFWDL ����WAIT�JN録��pnܷt�	TIMn����VAnp��_�UNITI�yL]Cg TRYn�u�dpMON_AL�IAS ?e	�phe5���� ��//'/9/�]/ o/�/�/�/P/�/�/�/ �/?�/5?G?Y?k?}? (?�?�?�?�?�?�?O O1OCO�?gOyO�O�O �OZO�O�O�O	__�O ?_Q_c_u_�_2_�_�_ �_�_�_oo)o;oMo �_qo�o�o�o�odo�o �o%�oI[m *������ �!�3�E�W��{��� ����Ïn������ /�ڏS�e�w���4��� ��џ������+�=� O�a����������ͯ x����'�ү8�]� o�����>���ɿۿ� ����#�5�G�Y�k�� �ϡϳ����ς���� �1���U�g�yߋߝ� H���������	��-� ?�Q�c�u� ���� ��z�����)�;��� _�q�������R����� ����7I[m *������ !3E�i{������$SMO�N_DEFPRO�G &����� &�*SYSTEM*��� $JO��RECALL �?}� ( ��}2xcopy �fr:\*.* �virt:\tm�pback@!=>�10.109.3�.132:598�4 e"n/�/�/�-}37%a?/Q/c$k/�/�? ?� 78$s:o�rderfil.dat�,�/�/~?�?��?}.8"mdb:�/[?4 f?�?	OO �%6/�/Z/�?}O�O�O �/EOWO�/�O__2? D?�?�?y_�_�_�?�? ]_f_�_	oo.O�O�O dOuo�o�o�O�OOo�O �o*_<_�_`_q ���_�_U�_�� �&o8o�o\o#���� $��oG��ol����!� 4F�j�{������ M��h�����0�Ï Տf�w�������?�Q� �����,�>�ǟb� s���������W���� ��(�:�ͯ^�oρ� �Ϧ���I�ܯ����� ��6�H�ѿ��}ߏߡ� ��O�ؿj�����2� ����h�y����A� S�����	��.�@��� d�u������߾�Y��� ��*�<���`�q �����K��� &�8�J��#� $��Q��l�/!/ 4���{/�/�/� C/U/��/??0B ��w?�?�?��/[? ��?OO,/>/�/b/ sO�O�O�/�/MO�/�O __(?:?�?^?o_�_ �_�?�?S_�?�_�_o�#n�$SNPX_�ASG 2����Ba�o  01Q%�#o�jo  ?�3fPA�RAM Be�La �	XkP�md1Pmh�d��C`5`OFT_K�B_CFG  �mcHe2cOPIN_�SIM  Bk��b);Es5`R�VNORDY_DOO  �e�eWr�QSTP_DSB�~�b�*kSR �Bi � &Ƚj��w�t�cTO�P_ON_ERR�d3b	�PTN �Be<��A�&�RING_PR�M�vrVCNT_�GP 2Be�aO`x 	���1P��������.gVDk�RGP 1v�a�`ҁ Bqď�.�@�R�d��� ��������П���� �*�Q�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ݿڿ����"�4�F� X�j�|ϣϠϲ����� ������0�B�i�f� xߊߜ߮��������� �/�,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZ�~���� ��� GDV hz������ /
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�?��?�?�?�?�?��PRG_COUNT�fs�<�IENBQ��EMAC�dNO_UP�D 1�{T  
O0R�O�O�O�O �O�O_-_(_:_L_u_ p_�_�_�_�_�_�_o  oo$oMoHoZolo�o �o�o�o�o�o�o�o%  2Dmhz�� �����
��E� @�R�d���������Տ Џ����*�<�e� `�r���������̟�� ���=�8�J�\��� ������ͯȯگ�� �"�4�]�X�j�|��� ����Ŀ�����5��0�B�L_INFO� 1�El@��	 eϩϔ���ϸ�@9�@??k�<��>�Ϻ���/HiB9�����{��H��bB/Hl������ A�����K� C�����
B���>�3���}�pz���\����C��F���������=�	Y=�J@YSDEBUG&@ʇ@�\�doI��SP�_PASS&EB�?��LOG ����A  \��K�b�  �kA\�?UD1:\��i���_MPC�݆EW�$i�A�� �A7�?SAV ��5A��������S�V.�TEM_TI_ME 1���@ 0�Ш���������MEMBK  �EkA����k��}�(�X|l@� @����Я�����Ȩ�	%
�� ��@
�L^p��〚����� �,>Pbt�����<e��/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"?4?F?��SKB�G�1A`V��?�?�?��7\�eFI2���9A�>A J��&O3I('!�;kO�:�O���N��` ��O�H0 �O_#_G_C�l_ ~_�_�_�_\�$�_�_ �oo%o7oIo[omo o�o�o�o�o�o�o�o�!3EWK?T1�SVGUNSPD��� '���zp2�MODE_LIMG ���vt2�p�qI���uuASK_OPTION��tJ����q_DI��?ENB  �5��� �BC2_GRP 2i5��	�A����9PCY@X�n|BCC�FG /��� 1�梏��`��*� �Ώ���=�(�a� L���p�������ߟʟ ��'��K�6�[��� l�����ɯ���د�#�+��=��p��� ��_�����ܿǿ ώ�  �L���(�N�<�r�`� �τϺϨ�������� �8�&�\�J߀�nߐ� �ߤ���������"�� 2�4�F�|�b�M���� ������b�����>� ,�b�t���T������� ������L: p^������ � 6$ZHj l~������/  /2/D/�h/V/x/�/ �/�/�/�/�/
?�/.? ?R?@?b?d?v?�?�? �?�?�?�?OO(ONO <OrO`O�O�O�O�O�O �O�O__8_�P_b_ �_�_�_"_�_�_�_�_ �_"o4oFoojoXo�o |o�o�o�o�o�o�o 0TBxf�� �������*� ,�>�t�b���N_�� ������(��8�^� L�������t�ʟ��� ܟ� �"�$�6�l�Z� ��~�����دƯ�� ��2� �V�D�z�h��� ����Կ¿�����"� @�R�d�⿈�vϘϾ� ���������*��N� <�r�`߂߄ߖ��ߺ� ������8�&�H�n� \����������� ����4�"�X��p��� ������B������� BTf4�x� ������, P>tb���� ���//:/(/J/ L/^/�/�/�/n��/�/  ??$?�/H?6?X?~?�l?�?�6�0�$TB�CSG_GRP �2�5��  ��1 
 ?�  �?�?�? !OOEO/OAO{OeO�O�K�2�3�<d�@ ��A?�1	 �HBL�H�0�F�DB$  C��2_&X��O_Cz&_n]A���H333?&ffo?���EA�_t�_~P �H���V̙U�PDH�_�]@���P�E�Qe�DaD" �A9oo�_(o�oLjX �FX�e�o�o�o�o@�o�o:Wf{<x�q	V3.00�2�	lr2dfs	�*�p�t�2�p �q<y �p�}��  �#�2��1J�2�3�=�qd�A�C�FG  �5��1 �0h����r�h������ ��0���;�&� _�J���n�������ݟ ȟ��%��I�4�Y� �j�����ǯ���֯ ����E�0�i�T��� ���2� ����οx�� ��7�"�[�F��j� �ϵ����ϔ�����!� �1�W��1�?|߈?�� �ߠ����������� B�0�R�x�f����� �����������>�,� b�P���t��������� ����(:�/Rd �������  "HZl*| ~�����/ / �D/2/h/V/x/z/�/ �/�/�/�/
?�/.?? >?d?R?�?v?�?�?�? �?�?�?�?*OONO<O rO`O�O�O�O�Ov�O �O_�O8_&_H_J_\_ �_�_�_�_�_�_�_o �_4o"oXoFoho�o�o �olo�o�o�o�o0 TBdfx�� ������*�P� >�t�b���������̏ Ώ����:�(�^�p� _����X�V�ܟʟ � �$��4�6�H�~��� ��`���دƯ��� � 2�D�V��z�h����� ��Կ¿����
�@� .�P�R�dϚψϾϬ� ��������<�*�`� N߄�rߨߖ߸ߺ��� �|��,�>���n�\� ~����������� "�4�F��j�X���|� ������������ B0fT�x�� ����,< >P�t���� ��/(//L/:/p/ ^/�/�/P�/�/V�/ ? ?6?$?Z?H?j?�? ~?�?�?�?�?�?O�? 2O OVOhOzO�OFO�O �O�O�O�O
_�O.__ R_@_v_d_�_�_�_�_ �_�_�_oo(o*o<o ro`o�o�o�o�o�o�o �o8�/�/bt L������ "��F�X�j�|�:��� ������ď����0� �T�B�x�f������� ���������>�,� b�P�r���������� ί����(�^�L� ��p�����ʿܿ��� ��¿H�6�l�Z�|� ~ϐ��ϴ������ ߀��D�2�h�Vߌ�v� s �ж� ����߶��$TBJO�P_GRP 2!�~�� / ?���	�����#������@� �0�  � �� � � �=�� @���	 �BL  f�?Cр D������[����<��B$\����@���?�33C�p���~�����f�x�x���*�;�2�������@��?�� �zX���s�A���� � ��S�Ʋ�>������;���pAW�?�ff�@&ff?�ff����~� �����x;7I
:v,�c?L������DH$ x{ ��@�33��"4�>������8�����Z�O�D"�#����xZVh9��� �������� �/=//�\/v/`/ n/�/�/�/b/�/?�/0�/,?]?��C���O���	V3.0~9�	lr2d�*�0�Ѷ?�7� E8� EJ�� E\� En�@ E�E�� �E�� E�� �E�� E�h �E�H E�0 �E� E��0��� E��0� �E�x E�X �F��2D�  �D�` E�0�P E�0$�00�@;�0G�0R@^op Ek�0u��0�@�0@�(�0� �E��0��0�X O9�IRzAF<�E��*�ߦO�B���CV����O��ESTPARS�@�������HRPABLE �1$���@��D�H�G *��I�G�H��H�׽��G	�H
��H�HKU���H��H�H�A+SRDI3_��J_\_n_�_�_�UdOo&k0oBoToHfoxn,RSo�� �Z 9K]o���� �����#�5�G� Y�k�}�����p�� IWЉ�o�o�o�o�_�_��_�_�_�X,R��NUoM  ~���B��� �@�@,R_CFG %���L�Z�@��IMEBF_TTQG���$P��VER�C�����R 1&;[ �8�?����T� ��ۏ  <�N�`�r� ��������̯ޯ�� �&�8�J�\�n���ɿ ������ڿ���"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�x��ߜ߮����� ������,�>�P�RR$�_���@�PMI_CHAN�� � ��DBGL�V����Q��E�THERAD ?UU���@d��b�*�<�X��ROUmT�!�j!p����a�SNMASK����255.����3�������3PO�OLOFS_DI�P����ORQC?TRL '+��c�OlT[���� ��� 2DV hz����Z���/SPE_DE�TAI��1
PGL�_CONFIG �-������/�cell/$CID$/grp1/@�/�/�/�/�/c�W� �/??*?<?N?�/r? �?�?�?�?�?[?�?O O&O8OJO�?�?�O�O �O�O�O�OiO�O_"_ 4_F_X_�O|_�_�_�_ �_�_e_w_oo0oBoTofoڎ}�_�o�o�o��o�o�od���m� �_Sew����_ �����+��O� a�s���������J�ߏ ���'�9�ȏ]�o� ��������F�۟��� �#�5�G�֟k�}��� ����ůT������ 1�C�үg�y������� ��ӿb���	��-�?� Q��uχϙϫϽ��� ^�����)�;�M�_��Z �User� View o)}�}1234567890�ߢߴ�����`����{�O#���v�2����T�f�x�������}�37����� �2�D�V���w�%�4 �����������
i�+%�5��dv�� ���%�6S *<N`r��%�7���//&/�G/%�8��/�/�/��/�/�/9/�/2 �lCamera��w/@?R?d?v?�?�?xbE3?�?�?�> ��OO&O8OJO\OR	  66�/?�O�O�O �O�O_�?*_<_N_�O�r_�_�_�_�_�_�/� 6��c_o*o<oNo`o ro_�o�o�oo�o�o &8�_�W���o �������o� �&�qJ�\�n����� ��K�WxK=���� (�:�L��p�����ߏ ��ʟܟ� ����5 ��\�n��������� ]�گ���I�"�4�F� X�j�|�#��W��ȿ ڿ����"�ɯF�X� jϵ��Ϡϲ������� ���Wn)�4�F�X�j� |ߎ�5ϲ�����!��߀��0�B�T����9 �ߕ����������  �%�7���H�m����P������V*	50M� &8J\�� ��K����� "����!0#;�{� ����|�// hA/S/e/w/�/�/B 5�K2/�/�/??/? A?�e?w?�?�/�?�? �?�?�?O�/���[�? SOeOwO�O�O�OT?�O �O�O@O_+_=_O_a_ s_O,Eg{
_�_�_�_ �_oo�O=oOoao�_ �o�o�o�o�o�o�_,E Ӌvo+=Oas� ,o������ '�9�K��o,E?���� ����͏ߏ��'� 9���]�o���������^�  b���� 
��.�@�R�d�v���<����   ��ğ �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� �����������ﰬ�  
^�(  }�ڐ( 	 .� d�R��v������ ������*��N�<�r�:8�̪ ���� ����N���#5G Y`��������� ��%lI[ m������� 2/!/3/zW/i/{/ �/�/�/�
/�/�/? R//?A?S?e?w?�?�/ �?�?�??�?OO+O =OOO�?sO�O�O�?�O �O�O�O__\OnOK_ ]_o_�O�_�_�_�_�_ �_4_o#o5o|_Yoko }o�o�o�o�_�o�o�o Bo1CUgy�o �o����	�� -�?�Q��u������ ��Ϗ����^�;� M�_�����������˟ ݟ$�6��%�7�~�[� m����������ٯ� ��D�!�3�E�W�i�{� ¯����ÿ
�������/�Aψ�h�@  c�pςϔ�c�j�N����+frh:\�tpgl\rob�ots\lrm2�00id��_ma�te_��.xml P�����0�B�T�f�0xߊߜߌ������� ������%�7�I�[� m���ߢ������� ���!�3�E�W�i�{� ������������� /ASew��� �����+ =Oas���� ���//'/9/K/ ]/o/�/��/�/�/�/ �/�/?#?5?G?Y?k? }?�/�?�?�?�?�?�? OO1OCOUOgOyO�N:��� jϸ��<< �� ?��K�O�O�O�O_�O _L_2_d_�_h_z_�_ �_�_�_ o�_o6oo�.oPo~o����(��$TPGL_OUTPUT 0���`  �e�o�o�o	-? Qcu����� ����)�;�M�_��q��e�@��`2345678901�� ����̏ޏ�������� �1�C�U�g�y��}�@����ӟ�����}� )�;�M�_�q�	���� ��˯ݯ�����7� I�[�m�������ǿ ٿ�������3�E�W� i�{ύ�%ϛ������� ��ߣ��A�S�e�w� ��!�3߿�������� ��'�O�a�s��� /������������ ��K�]�o�������=� ��������#��1�Yk}��9�b $$mb{�� �	�-QCu g������/ �)//M/?/q/c/�/@�/�/�/�/�/?}�A�?-???Q?c?u?�=@�O�?�?�J ( 	 ?�?�?OO 9O'O]OKOmOoO�O�O �O�O�O�O�O#__3_ Y_G_}_k_�_�_�_�_��_�_�_ooCo���  <<�/ xo�o�`go�o�o�o�o �o��do*<�oHr L^����� �&�8��\�n��V� ��>���ڏ�Ə�"� ��
�X�j������z� ��֟4�F�����&� T�.�@���������ү l�������>�P��� X��� �r���ο��� �b��:�L��pς� \ϊϸ�Ϡ��� ߚ� $�6��"�l����Ϣ� ��N��������� �2� ��6�h��T���� ����D�������R� d�>������������ |���$N���� ��0���� r8J�6�Z�l��Zb)WG?L1.XML�?���$TPOFF_�LIM _`�0[a��&N_S]V   �4%*�P_MON 1�We'$�0�02�)STRTCHK' 2We%&?"�VTCOMPAT�:(�!)&VWVAR� 3Z-�(>$ K�/ �/�0m"�!_DEFPR�OG %�)%IRVISIU �U?,_DISPL�AY �./2INST_MSK  �<� k:INUSsER�/q4LCK�<��;QUICKMExT0�?/2SCRE@�We�"tpscq4�1!@&I%"7@�_;IST�*%)RA�CE_CFG U4Z)�$o 	4�
?��HHNL C25>:7`�A�+ 2 �O�O�O_"_4_F_X_�jZ�EITEM 2�6�K �%$1�23456789y0�_�U  =<�_x�_�_�S  !�_k0�_Jo3�_ko �_�o�oo�o)o;o _o�o/U�o�o�o �o	�7�	�� ?����A���� ��Ϗ3�ۏW�i�{��� M���q���珏��� �A��e�%�7���M� ����������ů� ��a�	�������#�ͯ y������տ9�K�]� �����S�e�ɿq�� ����#���G���}� /ߡϳ�|��ϗ��ϧ� ��S�C�U�g߁ߋ�� ��[����߷��-� ?��c��5�G���S� ������w���)����� _�����^��y�� ���7�m -�=cu��� !�E�/)/� M/���Y/q//�/ �/A/�/e/w/@?�/[? �/?�?�/�??+?�?ʀDS�B7�O�:�g  uR�: �APOG9
 ]O�OjO��O(JUD1:\��L��AR_GR�P 18�[� 	 @P0�O[��O1__U_C_y_g^� �P�_�ZsQ�O�_�_�_�U?�  o)ko Io7omo[o�oo�o�o �o�o�o�o3!WEg�	�5��~	CSCB 29K o��#�5��G�Y�k�}����<UT�ORIAL :�K�OڏGV_CONFIG ;M��AMO�O9��OUT?PUT <I*���E������� ��џ�����+�=� O�a�'�v��������� ѯ�����+�=�O� a�r���������Ϳ߿ ���'�9�K�]�n� �ϓϥϷ��������� �#�5�G�Y�k�|Ϗ� �߳����������� 1�C�U�g�xߋ��� ��������	��-�?� Q�c�t���������� ����);M_ q�������� %7I[m~ �������/ !/3/E/W/i/z�/�/ �/�/�/�/�/??/? A?S?e?w?�%�t��? �?�?�?�?O!O3OEO WOiO{O�O�/�O�O�O �O�O__/_A_S_e_ w_�_�O�_�_�_�_�_ oo+o=oOoaoso�o �o�_�o�o�o�o '9K]o���o ������#�5� G�Y�k�}������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϴ� ���������!�3�E��W�i�{ߍߟ߂8������ߺѩ��� �?�1�C�U�g�y�� ������������� -�?�Q�c�u������� ���������); M_q����� ��%7I[ m������ �!/3/E/W/i/{/ �/�/�/�/�/�/�/? //?A?S?e?w?�?�? �?�?�?�?�?O?+O =OOOaOsO�O�O�O�O �O�O�O_O'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o"_5oGoYoko }o�o�o�o�o�o�o�o o1CUgy� ������	����$TX_SCR�EEN 1=����М}���\�n��������� J��I�����,�>� P�Ǐُ��������Ο ��W��{�(�:�L�^� p��������ʯܯ�  ��$�����Z�l�~� ������+�ؿO����  �2�D�V�Ϳz��� ����������oρ�.� @�R�d�v߈��Ϭ�#� ��������*��N���$UALRM_�MSG ?8��E� F�z����� ����������.�4��e�X���|���a�SEoV  o����_�ECFG ?v8�B�  u�@�  A  w B�t
 �� "s8�BTfx����������G�RP 2@�� 0v	 ,Na��I_BBL_NO�TE A��T?��l"r=��$q aDEFP�ROk�%o� (�%IRVISIONOy%���� /�8/#/\/G/�/�/�}/�/�/�/XFKE�YDATA 1B<8�8p v;>?P?'?t?�?]:�,(�?�?t(POINT  ]�?��>  OOK T� 	O�?NDIRE�CTOO CHO�ICE�?FOTOUCHUPqOrO�O �O�O�O�O	___?_ &_c_u_\_�_�_�_�_��_�_^9��/f�rh/gui/w�hitehome.png�_<oNo`o�ro�o�fpoint'o�o�o�o�o ��f  elook �b�o@Rdv�|indirec�o�����
�~choic&c�J�\�n�耏���`ftouchup�ʏ܏�� ���dfarwrg�L�^�p����� ���ß՟����� ��A�S�e�w�����*� ��ѯ�������=� O�a�s�������8�Ϳ ߿���'϶�K�]� oρϓϥ�4������� ���#�5�e:�a�s� �ߗߩ߻�������� �'�9���]�o��� ���F��������#� 5�G���k�}������� ��T�����1C ��Uy����� b�	-?Q� u�����^� //)/;/M/_/��/ �/�/�/�/�/l/?? %?7?I?[?�/m?�?�? �?�?�?�?z?O!O3O�EOWOiOkvK�>`����O�O �M�O�O�O�F,�_(_ �_L_3_p_�_i_�_�_ �_�_�_ o�_$o6oo ZoAo~o�owo�o�o�o �o�o�o2Vh Gߌ������? 
��.�@�R�d�v�� ������Џ�􏃏� *�<�N�`�r������ ��̟ޟ����&�8� J�\�n��������ȯ گ�����"�4�F�X� j�|������Ŀֿ� ��ϛ�0�B�T�f�x� ��Ϯ���������� ߩ�>�P�b�t߆ߘ� '߼���������� :�L�^�p����} ������ ��$�+�H� Z�l�~�������C��� ���� 2��Vh z���?��� 
.@�dv� ���M��// */</�`/r/�/�/�/ �/�/[/�/??&?8? J?�/n?�?�?�?�?�? W?�?�?O"O4OFOXO �?|O�O�O�O�O�OeO �O__0_B_T_�Ox_��_�_�_�_�_�_����[������o!o3moUogoAf,S�oK�o�o�o�o �o�o:L3pW ������ �� $��H�/�l�~�e��� ��Ə؏����� �2� D�V�e_z������� ԟ�u�
��.�@�R� d�󟈯������Я� q���*�<�N�`�r� �������̿޿�� �&�8�J�\�n����� �϶��������ύ�"� 4�F�X�j�|�ߠ߲� �������߉��0�B� T�f�x�������� �������,�>�P�b� t�������������� �:L^p� �������  $�HZl~�� 1����/ /� D/V/h/z/�/�/�/?/ �/�/�/
??.?�/R? d?v?�?�?�?;?�?�? �?OO*O<O�?`OrO �O�O�O�OIO�O�O_ _&_8_�O\_n_�_�_ �_�_�_W_�_�_o"o 4oFo�_jo|o�o�o�o �oSo�o�o0B�T+ V{�+ �����}{���v,Ï���,� �P�b�I���m����� ����Ǐ����:�!� ^�p�W���{�����ܟ �՟���6�H�'l� ~�������Ư�o��� � �2�D�V��z��� ����¿Կc���
�� .�@�R��vψϚϬ� ������q���*�<� N�`��τߖߨߺ��� ��m���&�8�J�\� n��ߒ��������� {��"�4�F�X�j��� ���������������� 0BTfx� ������, >Pbt�]��� ���/(/:/L/ ^/p/�/�/#/�/�/�/ �/ ??�/6?H?Z?l? ~?�??�?�?�?�?�? O O�?DOVOhOzO�O �O-O�O�O�O�O
__ �O@_R_d_v_�_�_�_ ;_�_�_�_oo*o�_ No`oro�o�o�o7o�o �o�o&8�o\ n����E�� ��"�4��X�j�|��������ď�Ƌ}������@���5�G�!�,3� x�+�������ҟ���� ݟ�,��P�7�t��� m�����ί�ǯ�� (��L�^�E���i��� ���ܿ� ��$�6� E�Z�l�~ϐϢϴ��� U������ �2�D��� h�zߌߞ߰���Q��� ��
��.�@�R���v� �������_���� �*�<�N���r����� ��������m�& 8J\������ ��i�"4F Xj������ �w//0/B/T/f/ ��/�/�/�/�/�/�/ Ϳ?,?>?P?b?t?{/ �?�?�?�?�?�?O�? (O:OLO^OpO�OO�O �O�O�O�O _�O$_6_ H_Z_l_~_�__�_�_ �_�_�_o�_2oDoVo hozo�oo�o�o�o�o �o
�o@Rdv ��)����� ��<�N�`�r����� ��7�̏ޏ����&� ��J�\�n�������3� ȟڟ����"�4�0�6��0���_�q���[�������,��诛���0� B�)�f�M��������� �����ݿ��>�P� 7�t�[Ϙ�ϼ��ϵ� �����(�?L�^�p� �ߔߦߵ������� � �$�6���Z�l�~�� ���C�������� � 2���V�h�z������� ��Q�����
.@ ��dv����M ��*<N� r�����[� //&/8/J/�n/�/ �/�/�/�/�/i/�/? "?4?F?X?�/|?�?�? �?�?�?e?�?OO0O BOTOfO=ߊO�O�O�O �O�O�?__,_>_P_ b_t__�_�_�_�_�_ �_�_o(o:oLo^opo �_�o�o�o�o�o�o  �o$6HZl~ ������� � 2�D�V�h�z������ ԏ���
���.�@� R�d�v��������П �������<�N�`� r�����%���̯ޯ� ����8�J�\�n���h����{@���{@���Ͽ��˿�'��,�X�� |�cϠϲϙ��Ͻ��� ���0��T�f�Mߊ� q߮��ߧ�������� ,�>�%�b�I���wO ����������%�:� L�^�p�������5��� ���� $��HZ l~��1��� � 2�Vhz ���?���
/ /./�R/d/v/�/�/ �/�/M/�/�/??*? <?�/`?r?�?�?�?�? I?�?�?OO&O8OJO �?nO�O�O�O�O�OWO �O�O_"_4_F_�Oj_ |_�_�_�_�_�_���_ oo0oBoTo[_xo�o �o�o�o�o�oso ,>Pb�o��� ���o��(�:� L�^�p��������ʏ ܏�}��$�6�H�Z� l���������Ɵ؟� ���� �2�D�V�h�z� 	�����¯ԯ����� �.�@�R�d�v���� ����п���ϕ�*� <�N�`�rτ�ϨϺ�@���������P����P����?�Q�c�;߅ߗ�q�, ����{������"�	� F�-�j�|�c����� ��������0��T� ;�x�_����������� ���_,>Pbt ��Ϫ���� �:L^p�� #���� //� 6/H/Z/l/~/�/�/1/ �/�/�/�/? ?�/D? V?h?z?�?�?-?�?�? �?�?
OO.O�?ROdO vO�O�O�O;O�O�O�O __*_�ON_`_r_�_ �_�_�_I_�_�_oo &o8o�_\ono�o�o�o �oEo�o�o�o"4 Fj|���� �o����0�B�T� �x���������ҏa� ����,�>�P�ߏt� ��������Ο��o�� �(�:�L�^�ퟂ��� ����ʯܯk� ��$� 6�H�Z�l��������� ƿؿ�y�� �2�D� V�h����Ϟϰ����� ���χ��.�@�R�d� v�ߚ߬߾������� ���*�<�N�`�r���[p���[p���������������,��8���\�C� ����y����������� ��4F-jQ� ������ B)fxW�� �����/,/>/ P/b/t/�//�/�/�/ �/�/?�/(?:?L?^? p?�??�?�?�?�?�?  OO�?6OHOZOlO~O �OO�O�O�O�O�O_ �O2_D_V_h_z_�_�_ -_�_�_�_�_
oo�_ @oRodovo�o�o)o�o �o�o�o*�oN `r���7�� ���&��J�\�n� ���������ڏ��� �"�4�;�X�j�|��� ����ğS������ 0�B�џf�x������� ��O������,�>� P�߯t���������ο ]����(�:�L�ۿ pςϔϦϸ�����k�  ��$�6�H�Z���~� �ߢߴ�����g����  �2�D�V�h��ߌ�� ��������u�
��.� @�R�d������������������$UI_�INUSER  �����  �����_MENHIS�T 1C�  ( �" ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,14������)n�621 �*<N` l,290���$���'v7//�A/S/e/�-�e�dit�IRVISION/�/�/�/ �/��7?I?[?m?xp?�48,2r?0�?�?�?�?���?O@-O?OQOcOuO��	A i	O�O�O�O�O�O _ O$_6_H_Z_l_~__ �_�_�_�_�_�_�_�_ 2oDoVohozo�oo�o �o�o�o�o
�o.@ Rdv�)�� �����<�N�`� r������O�Ȍޏ�� ��&�)�J�\�n��� ����3�ȟڟ���� "�4�ßX�j�|����� ��A�֯�����0� ��T�f�x��������� O������,�>�Ϳ b�tφϘϪϼϧ��� ����(�:�L�O�p� �ߔߦ߸���Y��� � �$�6�H�Z���~�� �������g���� � 2�D�V���z������� ������u�
.@ Rd������� �����*<N` ru������ �&/8/J/\/n/�/ /�/�/�/�/�/�/�/ "?4?F?X?j?|??? �?�?�?�?�?O�?0O BOTOfOxO�OO�O�O��O�O�O_���$�UI_PANED�ATA 1E����>Q � 	�}c/f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10nP�_Pice=TP&�_lines=3�nPcolumns�=4nPfonvP4�&_page=d�oub_P1_�)�prim�_�_  }�_oo1oCoUogo )io�oto�o�o �o�o�o�o/A(�eL�������  _ ���RdQ_Dc_u^2�_�_�V2��Wdual]����_ ����Ώ�����(� �L�^�E���i����� ��ܟß ��$�6��Z��~�@S������ į֯���M����B� T�f�x��������ҿ ����ݿ�,��P�7� t�[ϘϪϑ��ϵ�����s ~�	�A�S�e� w߉ߛ��Ͽ�2����� ��+�=��a�s�Z� ��~���������� ��9�K�2�o�V����� �*�������#5 ��Y��}���� �>��1U gN�r���� �	///?/����u/ �/�/�/�/�/"/�/? x)?;?M?_?q?�?�/ �?�?�?�?�?O�?%O 7OO[OBOOfO�O�O �O�OL/^/�O!_3_E_ W_i_{_�O�_?�_�_ �_�_oo�_AoSo:o wo^o�o�o�o�o�o�o �o+O6s� �O
_������ h9��_]�o������� ���ɏ�ԏ���5� G�.�k�R�������ş����������y��)�b�t���������) P��T�Я��1�C� U�g�ί��r������� �̿	��-�?�&�c� JχϙπϽ�M��s�{��$UI_POSTYPE  �u�� 	 ��� ���QUICKMEN  ����#���REST�ORE 1F�u�  �	��V��ߧӕ�V�m���� ��$�6��� Z�l�~���E����� ��������-�?��� z���������e����� 
.@��dv� ��W����O *<N`��� ��o�//&/8/ ��W/i/��/�/�/ �/�/�/�/"?4?F?X? j??�?�?�?�?�?�/ �?�?Oy?BOTOfOxO �O-O�O�O�O�O�O_��O,_>_P_b_t_.�S�CRE>�?C��u1sc���u2�T3�T4�T5*�T6�T7�T8�Q�SwTAT��� R�<�u��USER�P�_��Tks�SBd3Bd4�Bd5Bd6Bd7Bd8�Ba��NDO_CFG G��9�8����PD�Q,i��None1�#`_INFO 1H�u5�`P�0%z_�o M��o DV9z �o�����
����@�'��aOFF?SET K���aM�S��_������ Ǐ����*�!�3�}� 7���{�������ß� ����U�S�W�E�z��
j���V�a�aWO_RK L�mX����ۯ�O�"`UFR?AME  ���f��aRTOL_AB�RT>��cV�ENB�_�P�GRP 1M���O�Cz  A������a��ſ׿�@����1�R�=�U���an�MSK  h���an�N;�%�i��%'���p�_EV�N^����f�Ƅb2�No�
 h�a�UEV^�!td�:\event_�user\��"�C�7'�|�PF���S�P �%�spot�weldW�!CA6��]�o߱P��!�� 6���)���j����� \��<�N���r���� ���3���W���J� ������n������� /����e��F�X�|���
��WfŠ2O-i��8�Yk G��}� ���/�2/D// h/z/U/�/�/�/�/�/��/
??�/-?R?d?��$VARS_CO�NFI�`Po� F�PS�k<CCRG�bSo����?TuUD8� BHA�YpG�1C�A��G�A?�)@���=����CAA �3MRv��2Yo�c��P	�`ڢ%1:� SC130EFG2 *�O�@T�T�Y��j��5P�a�+AA@CC��> ��H�O!�_@(_U_zAP_}_�E/��A�0i_�_�2 B����Q�2�T a_�_A_o�_Bo-ofo Qo�ouo�o�oo�o�o��o�o,�_Pb�5TCC�3Z��/A�y/��;Dw0GF|0�[�o��02345678901�0�r��qA�1����@��Eq�5B�P�B�p�FL@AA:�o=L�RtEj��Aڡ�B g�3EA�Q�D��pb��?����"� 4�/�M�S�e�w����� ����я����B� =�O�u�s�������ү ͟ߟ��,�'��b� ]����������ɯۯ������tMODE�ȏ4 �tRSL�T \�<C%" �����o����<��s�p��ϵC�tSELE�C��;��qD�IA�_WO1]�5�R� �,	�	�Q���y�G�P� ǐ�;�=�RTS�YNCSE(Ѻ9���1��WINURLg ?��s@��π����,�>�P�r5I�SIONTMOU8(�u��� �h�s�^Sۣ�Sۥ�P�q FR:�\j�\DATA\�V� �� M�C��LOG��  � UD1��EX����1' B@� �����G�abriel_Faria���?�c��,@7F� n6  ������2� -ƌ�>A �  CE�4����>��TRAIN�;B4��d��pCE��� #`�=���ԍ�VB_�{ ( q	UyU_q� ������p%7Ib�STAW�`�y�B�@�����q$��e�_GE�s�a�{�  �
�W��08"'HOMI}N�pbSۮ�U �ؠ�ƱƱKAC�w����%JMPERR� 2c�{
   Q���/r��3�/�/? ??(?:?L?^?t?�?��?�?�?��S_�R�E�pd�utLEXz$e[�1-e/�VMPHASE � !%qCܲxqO�FF��_ENB { <�$VP2��_fSۯ�@x]#
���A@�T����B{�?s33������Am�B�D�Aʼxq
� i�-���*_>�<r�#`O� �D�"�e�֟������u_�� @�e�A���<q�*��1���9��-�u�_WBj� �_�_��o=��_�Wa_Vo�_ -o�_�o�o �o�ooco�o;o0B qoc�oo���o� �%�I[�K� Y�k��������� �3�ُ��1�C�U�� ������ܟ��� y��E�?���~����� џƯ���Q����� -�s�h���������߯ ��;�ݿ��+�]��� -ϓ��Ϛ�ɿ��%��� ����5�*�Y�K�}�r� �ϳ��ϣ߱��������QTD_FILTuE� j!+ ��& �Ȃ�I�[�m�� ����������C�3� �*�<�N�`�r����������	)SHIFTMENU 1k�-<�<%�?�4�� U,>�bt� ���	��?�(uL	LIV�E/SNAPi?vsfliv4N��� ION �l@U��menu ��_$/6/�����C�lY���MO�Cm� N�zQWAIT�DINEND  aD%�Ai"�&OKsHN�/OUT�/�(S�/�)TIM�%��	<G�/+=�/N;�/.:��/.:?�(RELE�KAtK�(TMz;e$=��#_ACT�sH�'A�(_DATA nU(B%8/^O���BRDIS��>��$XVRW!o�.�$ZABC_�GRP 1pU]Q ,e�2fO���ZD6@CSCH�Y q?I�!���KIPV"r�K%�h�__q_��_�IMPCF_GW 1s�I� P0R�f��_�Y�Ct�IP=pS� 	�_$o�  <�  �?�  ���;�4��aѿB`���DIa4���QaC����
_B��>a�>a��C��?����� � \����?C�� -o?oQocouo�o�m:��	'ooNa� ���C��F����������=�	Y=�J ewx^x�a����@���o�o�o�b0�o��o�D�PY u:_v�_�CYLIND�v�[ �:� ,(  *ȏٍA�ŏ0��&�� ?\� n������ǟ���� ��@�!�3�E���i�� ꟟���ï�������n��B2w�G*A ��_V���;��7�����F��:ז��A����SPHERE 2x���]�9ϭ�2� o�Vϓ�ۯ�����W� �Ϟτ�5��Y�@߲� �ߡ�������J����߀��1�x�U�g�y�@ZZ�6 �e&