��  I��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����SBR_T  � | 	$SVM�TR_ID  $ROBOT9�$GRP_N{UM<AXISQX6K 6NFF3 �_PARAMF	�$�  ,�$MD SPD_L�IT�?&2*�  � �E�NB�$$CLA�SS  ���������� V�ERSION��  0�~�IRTUAL���'  1 �� T���	M-10iA/7����  ai�S8/4000 �40A��
H1� DSP1-S1���	P01.0�5W,  	�  ��P�CR � ��C�����0���{  ���lr9  ?3!M�����  H��  �"`���
/m�~��  X���Z 
!
!������ ! ��
 1�2�
��?�0���VH.�������&����
= j ����� ?����������g�s� � �����w���)�.����NB� � d ���c �8 �:?�~��'b:
�c/ �/�/�/?��!,?��f<?a?s?�?���1�0���>���'�����3&2%-���0��?��_?����?�?&���<N`r�2|2����P�����}�9}�� ���� �W9 GA$((VA#�  h$ 4�����<����*��"r�:+�i�J | ��R 7�V$��?��d���z/��"�&؜/�/�D�/�_�_ �_�_!?�_E?o o2o�Do 5;����;�����8��&_88� ��8����_��$|#lFo�o����?�PB2/5 A2�m3|3<ONI
΄ �  V@�o�������{����<��9"�b8 l��  ���� �&��3 �'NHNH% �����2-����>��q k�� �a��:+p= � 	+��� MV$͘o�k �< 2|!� ����� ��r�l�&�c9�	`t # (��"� ��jTqrYa��K�]� o����_�� oɏۏ�����#�5�G���@��oNbiS�0.5/6�kx4�|4�o}�ϓ �o�_�K���q�/t�H���9�DsFp 82P�������;|�B'���S@A�S���� �����$x���  �� B�G�s;�T@;�����%}T���2�X���!�rY��~���
	�� �#�5���Y���}��������ſ׿����:�\d�N��R���x5|����Ԛ��~��J �p�~�<<���_@� ��{��"� �*�<���# �~v��!�V$�%�B�F�s�X@��x�"e�D�%¯ԯ ���������@���� v�?�Q�c�u���綠���N@�4JI�6|6d�{@��_d�R�a��t���t�a�_SnҴ��
�-8��0�o��� ����Ͻ��� �v�� uV$�����U`� J��s���Ta���D�ԄߖА�rY �+r��� t������ � �$���#5G�Yk�
������x�ҍ�Ng�	�t���� / /2/D/V/h/z/�/ �/�/�/�/�/�/
??.?@?P<�P?t?�?�? �?�?�?�?�?OO(O 0C��FO����O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_o^?&o8oJo\o no�o�o�o�o�o�o6O hOZO#~O�OXj| �������� �0�B�T�f�x����� ��
o�������,� >�P�b�t������o�� ��*<N�(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ȏ������ƿؿ��� � �2�D�V�ҟğn� ����������
�� .�@�R�d�v߈ߚ߬� ����������* N�`�r������� �����^ϐς�K��� �π������������� ��"4FXj| �����2�� 0BTfx�� �����R�d�v� >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?��?�?�? �? OO$O6OHOZOlO ~O���O/"/4/�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRo�?vo�o�o�o �o�o�o�o*�O �O�Os�O�O��� ����&�8�J�\� n���������ȏڏ� ��Zo�4�F�X�j�|� ������ğ֟�D�  �z��f�x����� ����ү�����,� >�P�b�t��������� �����(�:�L� ^�pςϔϦ�"���� 8�J�\�$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�ֿ �����������
�� .�@�R������ϛ��� �������*< N`r����� ��&��8\ n������� �/l�5/(/������ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?@OO,O >OPObOtO�O�O�O�O �OJ/</�O`/r/�/L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�?�o�o�o�o  2DVhz�O _�O�_0_�
�� .�@�R�d�v������� ��Џ����*�<� N��o`���������̟ ޟ���&�8��]� P������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� h�0�B�T�f�xϊϜ� ����������r�d�� ������t߆ߘߪ߼� ��������(�:�L� ^�p�������&� �� ��$�6�H�Z�l� ~�������0�"���F� X� 2DVhz� ������
 .@Rdv��� ����//*/</ N/`/���/x/�� �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4O�XOjO|O �O�O�O�O�O�O�O_ _�/�/6_�/�/�/�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�oNO(:L ^p�����&_ X_J_�n_�_H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ���o��ԟ���
�� .�@�R�d�v������ ���,�>���*�<� N�`�r���������̿ ޿���&�8�J�\� ���ϒϤ϶������� ���"�4�F�¯��^� د������������ �0�B�T�f�x��� ������������v� >�P�b�t��������� ������N߀�r�;�� ��p������ � $6HZl ~����"��� / /2/D/V/h/z/�/ �/�/�/�/BTf .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O��O�O�O �O�O__&_8_J_\_ n_�/�/�_ ??$?�_ �_o"o4oFoXojo|o �o�o�o�o�o�o�o 0B�Ofx�� �������v_ �_�_c��_�_������ Ώ�����(�:�L� ^�p���������ʟܟ �J �$�6�H�Z�l� ~�������Ưد4��� �j�|���V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ���������*�<� N�`�r߄ߖ����� (�:�L��&�8�J�\� n����������� ���"�4�F�X�j��� �������������� 0B�����ߋ�� ������, >Pbt���� ���//r�(/L/ ^/p/�/�/�/�/�/�/ �/ ?\%??��� ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O0/�O
__ ._@_R_d_v_�_�_�_ �_:?,?�_P?b?t?<o No`oro�o�o�o�o�o �o�o&8J\ n���O���� ��"�4�F�X�j��_ �_�_��o o���� �0�B�T�f�x����� ����ҟ�����,� >��P�t��������� ί����(���M� @���̏ޏ����ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� X� �2�D�V�h�zߌ� �߰�������b�T��� x�����d�v���� ����������*�<� N�`�r���������� ����&8J\ n���� ���6� H�"4FXj| �������/ /0/B/T/f/��x/�/ �/�/�/�/�/??,? >?P?�u?h?�� �?�?�?OO(O:OLO ^OpO�O�O�O�O�O�O �O __$_�/H_Z_l_ ~_�_�_�_�_�_�_�_ o�?|?&o�?�?�?�o �o�o�o�o�o�o
 .@Rdv��� ���>_��*�<� N�`�r���������o Ho:o�^opo8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� �����į֯���� �0�B�T�f�x�ԏ�� ��
��.�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ��p߂ߔߦ߸����� �� ��$�6ﲿ��N� ȿڿ쿴��������� � �2�D�V�h�z��� ������������
f� .@Rdv��� ���>�p�b�+�� ��`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?��?�?2DV O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�/�_�_�_ �_�_�_oo(o:oLo ^o�?�?vo�?OO�o �o $6HZl ~������� � �2��_V�h�z��� ����ԏ���
�fo �o�oS��o�o������ ��П�����*�<� N�`�r���������̯ ޯ:���&�8�J�\� n���������ȿ$�� �Z�l�~�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t������� �*�<���(�:�L� ^�p������������� �� $6HZ�� ~�������  2�����{�� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/?b?<? N?`?r?�?�?�?�?�? �?�?LOO��� nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_ ?�_�_o o0oBoTofoxo�o�o �o*OO�o@OROdO, >Pbt���� �����(�:�L� ^�p����_����ʏ܏ � ��$�6�H�Z��o �o�o���o؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .���@�d�v������� ��п�����t�=� 0Ϫ���Ο�ϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� H��"�4�F�X�j�|� ��������R�D��� h�zό�T�f�x����� ����������, >Pbt���� ���(:L ^p������&� 8� //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?�h?�? �?�?�?�?�?�?
OO .O@O�eOXO��� �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oop?8oJo\o no�o�o�o�o�o�o�o �ozOlO�O�O�O| �������� �0�B�T�f�x����� ����ҏ.o����,� >�P�b�t������� 8*�N`(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�ڏ����ƿؿ��� � �2�D�V�h�ğ�� ����������
�� .�@�R�d�v߈ߚ߬� ����������*�<� ��`�r������� ������&��ϔ�>� �����Ϥ��������� ��"4FXj| �������V� 0BTfx�� ���.�`�R�/v� ��P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O��O�O"/4/F/ _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodo�?�o�o�o �o�o�o�o*< N�O�Of�O�O_� ����&�8�J�\� n���������ȏڏ� ���"�~oF�X�j�|� ������ğ֟���V �zC���x����� ����ү�����,� >�P�b�t��������� ο*����(�:�L� ^�pςϔϦϸ���� ��J�\�n�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� 述���������
�� .�@�R�d�v����ώ� ��,���*< N`r����� ��&8J�� n������� �/"/~�����k/�� ���/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?RO,O >OPObOtO�O�O�O�O �O�O</_�Or/�/�/ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�oO�o�o�o  2DVhz� �__�0_B_T_� .�@�R�d�v������� ��Џ����*�<� N�`�r��o������̟ ޟ���&�8�J�� ����� �ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �z�0�T�f�xϊϜ� �����������d�-�  ߚ������ߘߪ߼� ��������(�:�L� ^�p��������� 8� ��$�6�H�Z�l� ~���������B�4��� X�j�|�DVhz� ������
 .@Rdv���� ����//*/</ N/`/r/�� ���/ (�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFO�XO|O �O�O�O�O�O�O�O_ _0_�/U_H_�/�/�/ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o`O(:L ^p������ �j_\_��_�_�_l� ~�������Ə؏��� � �2�D�V�h�z��� �������
�� .�@�R�d�v������ (���>�P��*�<� N�`�r���������̿ ޿���&�8�J�\� n�ʟ�Ϥ϶������� ���"�4�F�Xߴ�}� p������������ �0�B�T�f�x��� ������������,� ��P�b�t��������� �������߄�. �ߺ��ߔ���� � $6HZl ~������F� / /2/D/V/h/z/�/ �/�/�/PB?f x@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O��O�O �O�O__&_8_J_\_�n_�_�%�$SBR�2 1 5�P� T0 �  @?7 �_�_�_ o o2oDoVohozo�o �o�o�o�o�Q�o�_  2DVhz�� ������o��o @�R�d�v��������� Џ����*��N� 1�r���������̟ޟ ���&�8�J�\�?� ��c�����ȯگ��� �"�4�F�X�j�|��� q�����ֿ����� 0�B�T�f�xϊϜϮ��ϣ�~�_�����!� 3�E�W�i�{ߍߟ߱� �����������(�:� L�^�p������� ���� �����H�Z� l�~������������� �� 2D(�:�z �������
 .@RdvZ� �����//*/ </N/`/r/�/�/�/� �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �/�?O"O4OFOXOjO |O�O�O�O�O�O�O�O _�?0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>o"_boto�o�o�o �o�o�o�o(: L^pTo���� �� ��$�6�H�Z� l�~������Ə؏� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����Я���؟�*� <�N�`�r��������� ̿޿���&�
�4� \�nπϒϤ϶����� �����"�4�F�X�<� |ߎߠ߲��������� ��0�B�T�f�x�� n߮����������� ,�>�P�b�t������� ��������(: L^p����� ����$6HZ l~������ �/ /D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?6/v?�?�? �?�?�?�?�?OO*O <ONO`OrOV?h?�O�O �O�O�O__&_8_J_ \_n_�_�_�_�O�O�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�_�o 0BTfx� ��������o ,�>�P�b�t������� ��Ώ�����(�:� �^�p���������ʟ ܟ� ��$�6�H�Z� l�P�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ��ϴ�����*� <�N�`�r߄ߖߨߺ� ���������&�8�J� \�n��������� �����"���X�j� |��������������� 0BT8�J�� ������ ,>Pbt�j� ����//(/:/ L/^/p/�/�/�/�/� �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �/O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _ O@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo2_ro�o�o�o�o �o�o�o&8J \n�do���� ���"�4�F�X�j� |��������֏��� ��0�B�T�f�x��� ������ҟ��ȏ�� ,�>�P�b�t������� ��ί������:� L�^�p���������ʿ ܿ� ��$�6��D� l�~ϐϢϴ������� ��� �2�D�V�h�L� �ߞ߰���������
� �.�@�R�d�v��� ~߾���������*� <�N�`�r��������� ������&8J \n������ ����"4FXj |������� //0/T/f/x/�/ �/�/�/�/�/�/?? ,?>?P?b?F/�?�?�? �?�?�?�?OO(O:O LO^OpO�Of?x?�O�O �O�O __$_6_H_Z_ l_~_�_�_�_�O�O�_ �_o o2oDoVohozo �o�o�o�o�o�o�_�o .@Rdv�� ��������o <�N�`�r��������� ̏ޏ����&�8�J� .�n���������ȟڟ ����"�4�F�X�j� |�`�����į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ������Ŀ��(�:� L�^�p߂ߔߦ߸��� ���� ����6�H�Z� l�~���������� ��� �2��(�h�z� ��������������
 .@RdH�Z�� �����* <N`r��z� ���//&/8/J/ \/n/�/�/�/�/�/� �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? �/O0OBOTOfOxO�O �O�O�O�O�O�O__ ,_OP_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^oB_�o�o�o�o�o �o�o $6HZ l~�to���� �� �2�D�V�h�z� ����������
� �.�@�R�d�v����� ����П�Ə؏�*� <�N�`�r��������� ̯ޯ�����
�J� \�n���������ȿڿ ����"�4�F�*�T� |ώϠϲ��������� ��0�B�T�f�x�\� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ ���2DVhz �������
/ /./@/$d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?V/�?�?�? �?�?�?OO&O8OJO \OnO�O�Ov?�?�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�O�O�_ oo0oBoTofoxo�o �o�o�o�o�o�o�_ ,>Pbt��� ������(� L�^�p���������ʏ ܏� ��$�6�H�Z� l�