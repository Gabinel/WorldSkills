��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� � P�COUPLE,  o $�!PPV1OCES0�!H1�!��PR0�2	 � $SOFT��T_IDBTOT_AL_EQ� Q1�]@NO`BU SPI�_INDE]uEX�BSCREEN_��4BSIG�0�O%KW@PK_F�I0	$TH{KY�GPANEhD� � DUMMYE1d�D�!U4 Q_���ARG1R��
 � $TIT1d ��� 7Td�7T� 7TP7T55V6�5V75V85V95W0 5W>W�A7URWQ7UfWU1pW1zW1�W1�W� 6P!SBN_CmF�!�0$!�J� ; 
2�1_CM�NT�$FLAsGS]�CHE"{$Nb_OPT�3��(CELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1�UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t��d�MO� �sE' � [M�s���2�REV�BI�LF��1XI� %�R�  � OD�}`j�$NO`M�+��b�x�/�"u�� ����Q�X�@Dd p =E RD_Eb��?$FSSB�&W`�KBD_SE2uAUG� G�2 "_��B�� V�t:5`ׁ8QC �a_EDu �� � C2�2�`S�p�4%$l �tO$OP�@QB�q�y�_OK���0, P_C� y��dh�U �`/LACI�!�a��x�� FqCOMM� �0$D��ϑ�@�p�X��ORB�IGALwLOW� (KtD2�2�@VAR5�0d!�AB e`BL[@S � ,KJqM�H`9S�pZ@M_O]z�ޗ�CFd �X�0GR@��M�NFLI���;@UIRE�84�"� �SWIT=$/0_NZo`S�"CFd0M�� �#PEED��!�%`���p3`%J3tV�&$E�.�.p`L��ELBOF� �m��m�p/0$��CP�� F�B�����1��r@1J1E-_y_T>!Բ�`���g���G� }�0WARNMxp��d�%`�V`NST�� COR-rF�LTR�TRAT� T�`� $AC�CqM�� R�r$�ORI�.&ӧRT��SFg CHG*V0I�p�T��PA*�I{�T�P�|�� � �#8@a���HDR�B�ą2�BJ; �C��3��4�5�6�7
�8�9�4��x@�2� @� TRQB��$%f��ր���֣_U���ѡ�Oc <� ����Ȩ3��2��LLECM�>-�MULTIV4�"�$��A
2q�CHILaD>�
1��z@T_1b�  4� STAY2�b4�=@�)2�4����@�� | 9$��T�A�I`�LE��eTO���E��EXT���ᗑ�B�᎞22�0>���@��1b.'��}!�A�K�  �"K�/%��a��R���?s  =�O�!M��;A�֗�qM�� 	�  =��I�" L�0[��� R�pA��$JO�BB������TRIGI�# dӀ���� R�-'r��A�ҧ��s_M��b$ tӀ3FL6�BNG�A��TBA� ϑ�!��
 /1�À�0���R0�aP/p ����%��|��Bq@W�
2J�W�_RH�CZJ�Z�_zJ?�D/5C@�	�ӧ��@��Rd&������ȯ�q�GӨg@NHANC��$LG/��a2qӐ� ـ@��A�p� ���aR��>$x��?#3DB�?#RA�c?#AZt@�(.�����`gFCT����_F�L�`�SM��!I�+ lA�%` �` ���$ /�/����[�a���M�0\��`��أHK���AEs@͐�!�"WꍠN� SbXYZ�W�`�"����6	�������'  E. II��2�(p�STD_C�t�1Q���USTڒU�)�#�0U[�%?IO1��� _Up�q��* \��=�#AOR@zs8Bp;�]��`O6  RSY�G�0�q^E�Up��H`G�� ��]�DBPXWORK��+* $SKP_��p��A�TR�p , �=�`����Z m�OD3��a _�C"�;b�C� �GPL :c�a�tőS�D�W�3Bb����P�6�P )DB�!�Y-�B APR��
I�8Ja3��. /�u�\������LuY/�_�����0�_����PC�1�_����~�EG�]� 2��_�SVPRE.��R3�H $C��7.$L8c/$uSނ�z IkINE�WA_D1%�ROyp��ŀ����q�c7 t@�fP�A���RETUR�N�b�MMR"U���I�CRg`EWM�@�SIGNZ�A� ���e� 0{$P'�1$P� &m�2p�p'tm�+pD�@ �'�bdNa|)r�GO_AW ���@ؑB1I�CYSd�(�CYI�4��B�`1w�qu��t2�z2�vN�}��E}s�DEVIs` 5� P $��RB���I�wPk��IG_BY���"�T7Q��tHNDG�Q6� H4��1�w��$DSBLC��o��vhg@��|tL��7O��f@]���FB���FEra8�ׂ�t}s����8> i�T1?���MCS���fD �ւ[2H� W��EE���%�F����t����9 Tx�p��x�NK_N:�Ԅ���U��L�wHA�vZ' ~�2���P�~r�q7: �=MDLn��9�ጂٱ h����!e����J��~�+����,�N�D����3��ՒG!a�qSLAd�7;  ��INP��"������}q_ �4<�0�6`C� NU�� � D�Lק��SH!�7=M��q���ܢӢ���g���?>P +$ٰ��٢��^��^�Y�FI B\��Ă��'A�	'AWl�NTV���]�V~�X�SKI�#T���a�ۺ�T1�J�3:3_�P�SAqFN���_SV��EXCLU��N@J�DV@L��@�Y��<��S�HI_V
0\2�PPLYPRo�HqIM�T�n�_MLX�}�pVRFY_�C:l�M��IOC�UCC_� ����O�Fq�LS�0v�FT4QI�����@P�E�$�t��A��CNF�t�6եu��pm�4AC�HD�o������AMFC CPlV�TQpTP?�� �� ?`Ɵ@TA�@�0L@ ���N��]� @$����T��T! S���x�te@{RA DO��� w2���!In��_1�#�H!�(̔�΀K��B�2��_MARGI�$����A ��_SG5NE�C;
$�` �a^aR0��3��@ B���B��ANNUN��P?���uCN@ �`%0����� ���B�EFc@I�RD @bQ�F���4OT�` �sFT�HR,Q��CQ0�-M��NI|RE������AW���DAY=CLOAD�t;T|��<S5}�EFF_A+XI��F`1QO3�O��Eq��@_RWTRQE�G���V�0RQ�2Evp ��|�F�0f�R0| �tM�AMP�}E<� H 0��`œ^�`Ds�DU��`���BCAr� �I?�`N ErIDLE_PWRIh\V!n0V�wV_[ ||�� �DIAG�5J� 1$V�`SE�3TQl�e�`�Pl�^E_��Y�VE� �0SWH�q(� �b|��Gn�OHxP�PHZ�IRAl�B �@�[��a�b�1� w3�O � ��v�|��I�0 �pRQD�W�MS-�%AXx{6Y�LIFE�@�&�MQy�NH!Q%H��F#C����CB0��mpN$�Y @�aF3LAl���OV0]&�HE��l�SUPPIO�@u�y��@_�$��!_X83�$gq�'Z�*W�*B1�'T�#�`�k2XZáY�Y2�D8CY`T@�`N����f� �C�I2ICTA�K =`�pCACH�ӫ�3����I��bNӰU7FFI� \��@���;T��<S6CQ.�M�SW�5L 8	�K�EYIMAG�cTMLa��*Ax�&E���B>��OCVIER-awM ��BGL��<��y�?� 	���j�4N�:�ST�!�BP�D,P�D�x�D��@EMAI��a��M�r�FAUL|RObB�c�� sp�UʰMA"`T'`E�P�< $S�S�[ � ITw�BUF��7y��7�tN[�LSUB1T�Cx�o�R�tRSAV|U>R'@c2�\�WT���P�T�*`Sn�_1PbU��F�YOT�bK��P��aM��d���WAX���2��X1P��S_G:H#
��YN_���Q <Q�D��0��U�M�� T�eF�`|�\�DI�ҏEDT_Pɰ:�R$��b�GRQM�&��Jq��a���׀��Fs� oS (�SVqp�B��4�_�.��a��T� �@���Bn�SC_R]1IK>B'r��$t��R"A#u�HN�aDSP:FrP�lyIM|Sas�qz��aB� U>w� <1%sM�@�IP��s��0`tT!Hb0ЃTr��T`assHS�cCsBSCʴq0� V�����S�{_D��CONVE�AG���b0^v1PFH�y�dCs�`&a?ASC8���sMERg��a�FBCMPg��`E�T[� UBFU&� DU%P�D�:1�2�CDWy�p�P�CGM�[@NO6�:�V� ��� ���P���C"�����w��A��|`��WH *�LƠ�Cc�W����Y� 賂��р�q�|�P��A��7}�8}��9}�H ���1��1���1��1��1ʚ1�ך1�1�2��2T����2��2��2��U2ʚ2ך2�2�3��3��3����3���3��3ʚ3ך3��3�4��QEX	T[�X[b�H``t&�``z�k`˷$���F{DR�YTP�V��RK"	��K"R�EM*F��]"OV�M:s/�A8�TRO�V8�DT�PX�MX�g�IN8ɉ W��INDv�H2
�ȕ`K ^`G1a�a��@Q%79Da�RIV��u"�]"GEAR:qIO.K(�H4N�`����,(�F@� I3Z_MsCM<0K! �F� 9UT���Z ,�TQO? b�y@t�.G?t�E |�p.�>Q����[ �5Pa� RI�E���UP2_ \ �@=STD	p<T�T���������a>RB;ACUb] T��>R
�d)�j%C�E��0��IFI��0��i�{��4�PTT��FLU=I�D^ �?0gHPUR�gQ�"�r�aP�4P+ I�$��]Sd�?x��J�`sCO�P�SVRT��>N�x$SHO* ��CASS��Qw%�pٴBG_%��3��࣓��FOR�C�B��o�DATAZ��_�BFU_�1�b:b�2�am=mm�b0���` |��NAVN	`������$��S�Bu#$VIS�I���2SC	dSE������V��O��$&�BK�� ���$PO��I���FMR2��a ��	��` #��&�8�O� �(�_����+IT_^�ۄ)M������DGCLF�DG�DY�LD����5�Y&��Q$Y�M됇Cb�N@{	 T�F9S�P�Dc P��W|�cK $EX_W�nW1%`]��"X3��5��G+�d� ���SWeUO>�DEBUG���-�GR��;@U�B�KU��O1R� _ PO_ )���t��M��LOOc>!SM� E�R�a���u _E e �>@�G�TERM�`%fi'�ORI�ae gi%y�SM_�`>Re hi%V�(�ii%3UP\Bjg� -���e���w#� f��G�*E�LTO�A�bF�FIG�2�a_���@�$��$g$UFR�b�$�1R0օ� OT_7F�TA�p q3wNST�`PAT�q<�0�2PTHJ�Ԁ�E�@�c3ART��P'5�Q�B�aREyL�:�aSHFT�r(�a�1�8_��R��уJ�& � $�'@i�p
����s@bSHI�0�Uy� �QAYLO�p�Oaq�����18����pERV��XA ��H��m7�`�2%�P���E3�P�RC���A�SYM�a��aWJ07����E�ӷ1�I��ׁUT�`Oa�5�F��5P�su@J�7FOR�`M  �O!k]��5&�0L0���sHOL ;l �s2XT����OC1!>E�$OP��q�n���$�����d$��PR^��aOU��3e��R�5e�X|�1 �e$PWR��3IMe�BR_�S�40�� �3�aUD���`t�Q�dm��$H�e�!�`ADDR˶HBR!G�2�a�a�a ���R��[�n H��S ����%��e3��e���eư�SE��L�HSv�MNu�o��`�Pªq��0OL�s�߰`ڵ�I ACR�O��&1��ND_C�s��AfdK�ROU	P��R_�В� �Q1|�=�s���y%��y -��x���y���y>�=�A��Ҁ�AVEDȻw-��um&sp3 $���P_D�� ���'rPRM_���HTTP_�H�[�q (ÀOBJ���b �$˶LE�~3�P��\�r � Q���ྰ_��TE#�ԂS�PIC��KRL~PiHITCOU�!��L���PԂ���0���PR��PSSB�{��JQUERY_F�LAvs�@_WEBwSOC���HW��#1��s�`<PIN'CPU(���O��� g�����d��t��O���IOLN�t� 8��R��$�SL!$INP7UT_U!$`���P  ֐SL.���u���2�.���C��B�IOa�F�_AS=v�$!L+ਇ+�A��bb�41�����Z@HY�ʷ����#qe�UOP:w `v�ϡ˶�� ��������"`PIC`����� �	�H�IP�_ME��v�x X�v�IP�`(�R�_N�p�d���Rʳp�ױQrSP �z�C��#BG(� ��M�Av�gy lv@CTApB��AL TI�3UfP�_ ۵�0PSڶBU_ ID� 
�L � ``�a�����0z)�"���ϴ�NN�_ �O��IRCA_C}Nf� { �Ɖm-�CYpEA�� ������IC�ǫ�tpxR�=QDAY_
��NTVA�����p!��5����SCAj@F��CL�
����
���v�|5�VĬ2b�l�N_�PCV�n�
���w�})�T��S������
��e���T� 2G| $� �v�~�8�֣�ذLAB1��\_ ��UNIX���� ITY裪��ea��R� ��<)���R�_URL���$A;qEN ���s`vs�TeqT_U���iJ��X�M�$���E�ᒐR祪�� A��,���JH���FL�y��= 
���
�wUJR|U� ���AF�6G��K7��D>��$J7�s��J8B*�7���3�E�7���&�8\�)�APHI�Q4�y�DkJ�7J8R��L_K�E'�  �K�͐LMX� � �<U�XRi�����WATCH_VAZqxu@AំFIEL`�b�cyn���:� � bu1VbwPCTX��j���LG~E��� !��?LG_SIZ΄�`[8Zm�ZFDeIYp1!gXb Z W �S`�8�m���� �b ��A�0_i0_CMc3#�*�'FQ1KW d(V(Bbpo  pm�p� |Io�`1 pb pW RS��ޜ0  (C�LN��R�۠�DE6E3����c�i��r�PL#�DAU"%�EAq�͐�T8". GqH�R��y�BOO�a?�� C��F��ITV�l$A0��RE���(SCRX�����D&�ǒ�qMARGI4�Sp�,����T�"$�y�S��x�W�$y��$��JGM7MN3CHt�y�FN��61K@7r�>9UFL87@nL8FWDL8HL�9STPL:VL8"�L8,s L8RS�9HOPh;��C9D�3R��}P�'IUh�`4�'�5$ d��S2G09�pPOWG��:�%�3,64��N9E]X��TUI>5I�  �ӌ�����C3�C<0'�,�o:��&�@�!9NaqvcANAy��Q��AI]�gt7Ӝ�D�CS���cRS�cRRO�XXOdWS�ÂRoXS{X�(IGNp 
Ђp=10 ��[TDEV�7�LL��Y"*�C �4	 8�Tr$f/�Л�����3A�a�B	 W�萦�Oqs�+S1Je2Je3Ja��8�BSPC � �ƋG`-T��%��Q�T��r@�&E�fST�R�9 YBr�a �$E�fC�k�g��fp	v9�CB� L�� ��� ��u�xs뀔�g��q�jt��!�#_ ���ʐv�#Ӡ �s� �MC�� =���CLDP᠜�TRQLI ���y�tFL���rQ��s5�1D���w~�LD�u�t�uORG���1�?RESERV��M�ຓM�Œ�t��� �� 	�u�5�t�uS�V��p��	1���>��RCLMC��M��_�ωА��_C�M�DBGh�I�����$DEBUGMA�S������U�$T�8P��EF�d��pF�RQҤ� � �K	HRS_RU�4�bq��A��$EFgREQ6u!$0YOVER�k�t�f�PU1EFI�C%Gq�� �
Y��z�� \����E�s$U�`��?���
�PSI`��	��C A ��ʲ�σUY�%��?( 	��MI;SC�� d��akRQ��	��TB� �� ���A��AX��𑧪�EXCE�Sg�9d�M�H��9�u���}qd�SC>�` � H�х�_�����������p�KE��+�� &�B�_, FLICBtB�� QUIRE CMEOt�O��얩qLdpMD� �p{!���5b���$L�M#ND!��I�����L �D;
$INAsUT�!
$RSM�ȧPN���C����PSTLH� �4U�LOC�fRI�"��eEX��ANG�.R.���ODA]�Řq��� �RMF 0����icr�@mu�Ŝ�$�SUPiu��F�X��IGG! � ���cs�F�cs 
Fct��ޒ�b5��`E؀�`T�5�tC��g�T!I��7 ;��M���7� t�MD���A)��XP��ԁ��H��.���DIAa��Ӻ�AW�!��0af���D@#�)֡O�㥀��� -�CUp V	����.���O�!_��ᜃ �{`�c����	�� |�P|��0� ���P{�KEB��e-�$B��o�=pND2xւ����2_TXlt�XTRAXS����&��LO: ����&}�L���C�.��&�[�RR2h���� -�!A�� d$CALI����GFQj�2F`RI�Nbn�<$Rx�S�W0ۄ���ABC��D_J��{�q���_J3��
��1S�P, �q�P����3P��H�9pq�#J�h3n���O�QIM���CSKP�zb7$?SbJ+ᯂQb�py����_AZ���/�EL�Q.ցO�CMP�ð�� R1TE�� �1�0 �F��1��@ Z�SMG�0�Э�JGΊpSCLʠ��SPH_�P��f��q�=u�RTER��n�IPk�_EP�q�`aA� �c���DI��Q23UdDF � ���LW�VE�L�qINxr�@�_�BLXP.��Y/�J`��'$"pIN����]�C�9%�".�t8!6p_T� �F% a"���^$��k)�F~pDHʠ��\�9`�$Vw��_�Aa$=��~�&A$���S�h��H �$BEL� m���_ACCE� x	8�0IRC_��q�@�NT��c�$PSʠ�rL� ��M4�s9 .7��GP/6 ��9�7$3�73S2T�͡_Ga�"�0�1��8�n1_MG}�DD�1�~�FW�p��3�5�$32�8DEKPP�ABN[7ROgEE�2KaBO�p�Ka���1�$USE�_v�SP��CTR�TY4@� �� <qYNg�A�@�FR �ѢA!M:�N�=R�0O�v1�DINC(��B�4p���GY��ENC��L��.�K12��H0I�N�bIS28U��ON�T�%NT23_�~�fSLO�~�|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1�����PERCH  �S��� �W���Sl� �R��l����E�0�0PAS2EeL�DP7��ONUЉZ�f�VTRK�RqAY"�?c� �aS2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gB�T�DUX �2S_BCKLSH_CS2 Fu:��V���C-�esR�oz�A�CLALM�JT@��`� �uCHK�e ����GLRTY@pн�8T��5���_��N�T_UM3��vC3�p�1Z���LMT���_LG��%���0�E *�K�=�)�@5F�@8 09�Nb��)hPC�Q)h�HТ��5�uCMC����0�7CN_��N����;SF�!iV �B��.W���S2/�Ĉ7CAT�~SH�Å� �4 V�q/q/V�T1���0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e�0�R� @B�_Wu�d��!a��#`��#`�I*h�Iv�I�#F��S��:��I�0VC00��֢1ܮ�0��JRKܬ!��<�KDBXMt�<�M��_DL�!_bGRV�g�`��#`��#A�H_p%�?��0��COS��� ��LN#���ߥŴ � ��=������꼰�b<�Z���VA�MYǱ�:ȧ��᯻[�THE{T0�UNK23�#؅��#ȰCB��CB�#Cz�AS�ѯ�0���#����SB�#��N��GTSkZAC�������&���$DU�phg6�j��E��%Q%a_��x�NE
hs1K�t�� y�A}Ŧկ׍������LPH����^U��S ߥ����������!�(�(Ʀ�V��V�غ ���V��V��V
�V��V&�V4�VB�H���������d�����H�
�H�H&�H4�H*B�O��O��Os���UO��O��O
�O�UO&�O4�O(�F����	���SPBALANCE_J��6LE��H_}�S�P>!۶^�^��PFULCb�q����K*1�UTOy_�p�uT1T2�	
22N�q2VP�M@�a� i�Z23	qTu`�O�1Q�INSE9G2�QREV�P�GQDIF�ep)1�lU�1��`OBK�qj�w2,�VP�qI�?LCHWAR4B�B�AB��u$ME�CH��J��A��vAX�aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ֯@�C1_ɒT �� x $W�EIGH�@�`$ȹ�\#��I�A�PIF�vA�0LAG�B��S��B:�BBIL�%O1D�`�Ps"ST0s"P:�pt � N�C!
L �P 
P2�Aɑ�  2��Tx&DEKBU�#L|0�"5�OMMY9C59N���$4�`$D|1 aq$0ېl� > �DO_:0AK!� �<_ �&� �q�A��B$�"� NJS�8_�P�@� �"O�p �� %�T7P?Q��TL4F0TICK,�#�T1N0%�3=pB�0N�P� u3�PR\p��A��5��5U0PR�OMP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a��@RU�COD�#F9U�@�&ID_�P�E�82B> G_SUFF�� �#�AXA�2DO�7/�5� �6GR�#��DC�D ��E��E-��DU4� u�_ H_FI�!�9GSORD�! R 236s�HR�A>N0$ZDT�E=!|� X5�4 *WL_NA�1�0�R�5DEF_I�X�RF �T�5�"�6�$�6�S�5�UFISm�#�m1|Ј�40c�3�T6�44􁆂�"D� ?rfd�#�D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D�S �D�U�D>b�B�c�E�S �Dd�B�&2v2a�C� ʑ�E�R�E�S�C9wwu�H�0P} d�0,a�ТF0W�h�u�c=!T�E�qY4� >�!LOMB_�r�w�0s"VIS��IT�Ys"AۑO�#A_�FRI��~SI,a�n�R�07��07�)3�#s"W�W�Q���%�_���AEAS {#�B��|�x`WB8��45�55�6|#OR�MULA_I����G�W� h �
>75COEFF�_O�1&)��1��Gdo�{#S� 52CA� �:?L3�!GRm� ?� � $�`�v2X�0TM�g���e��2�c��3ERIT��d�T� �  �L�L�Dp`S��_SVLkd��$�v� �.����� � ��SE;TU,cMEAG@�@�Πt �!HRL � �3 (�  0��@l��l��aw��R�0$�a�a}d]�d��B��Ay`Gax`��[�:�k@REC[Qq���QSK_A y��� P_!1_USER�����*���VEL����-��!��IzPB�MT�1CFG��� � �0]O�NO#REJ �0l���[�?� 4 e���"�XYZ<SB� x3:!��_ERRK!C� U ѐ�1�@c��Ȱ�!�>�B0BUFINDX���P� wMORy�� H_ CUȱ�1��dAyQx?�I>Q$ �+�a����� \�G�{�� � $S�I�h��@2	�VOxv�q�- OBJE| w�ADJUF2yĈ��AY�����D��O�UKP����AMR=�T��-���X2DIR����Xf�1�  DYNt�0�-�T�� ��R��0� ����OPWOR�� ��,B0SYSB9U����SOPo��$�z�Uy�XP�`K���PA�q������+OP�@U���}x�"1��IMAG۱1_ �п"IM.����IN������RGO�VRD"ё�	���P ����  >gplcC���L�`BŰ?l�PMGC_E�P�1N��Mr�1212R�"�sSL| ��� �R �OVSL=S�rD#EX\a`��2�:�_"���P#���P ������2�C �P�>���#�_ZER�l���:���� @h��:��O�@RIy��
[�g@e���s�P��PL���  _$FREEY�EU�Q~�Z��L����yT�� ATUSk��,1C_T�����B ������p�Vc1��P��� Dc1�к���LQ����MQ��ۡL�XE��x�5IP�1�W�` ��UP��H`�&aPX;@��43�����PGY��>g�$SUB����q���JMPWA�IT~ ���LOWp���1wē CVF_A��0��R�Z��C�C �R$��28IG�NR_PL��DB�TB� P*a�BW�@.t�U�0-IG���!@I�TNLND,�RBѡb�N!@���PEED~ ��HADOW� ��t����E������PSP]D��� L_ A��0�P���	#UNq �d �RP (�LYwP�a����PH_P�K���b�RETR#IE��x���2�R!vD@FI��� ���V �$ 2�d�D�BGLV<LOGgSIZz�baKT�U���$D��_T-XV�EM�Cڡ)��� �-R�#�r��CHECKz����L��%�ϰq)�L��NPA�`TJ"�����)1P����
�AR@�"�BC =Sa��O�@����ATTS�u���&� w�^a�3-#UX�^�4�PL�@Z��� $d��qSWIT�CH�h�W��ASr��f�3LLB���� $BAr�Dvc��BAMi�h�6I��(@J5���N�UB6[F
A_KN�OWK3qB"�U��A�D+Hc� D��IPAYLOAq�9p�C�_���GrѼGZ�CL�qAj��PLCL_6� !4��BOA�?�T7�VFYC�Ӑ�Jp��D�I�HR�Ր�G�TB��6�JL(�zQ_J�A �B�AND����T�BQ��q��PL@AL_ ��0 =�TAe��pC��D�CE���sJ3�P�V� T��PDCK^�)b��C}OM�_ALPH�S�cBE<�߁�_�\��X�x\� � ����OD_1�J2�DDM�AR<�h�ex�f�cQ�TIA4�iu5�i6��MOM(�@�c�c�c�c�cV�B� �AD�cv�cv�cPUBP�R�d<u�c<u��b}"�1���� L$PI$��pc���G�y��I�yI�{I�{I�s�`�A���v��v�J�b��a��HIG�3��� 0���5�0�f�?��5N�5�SAMP D Ƣ�0����;@�S ��с6���1� ��� ���`���`1�@K�P��`腽P�H��IN1��P��8�T��/��:�z�Q�z���G�AMM&�S���$GET�����D�^d>�
$�PIBRt��I��$HI��!_���1��E=��1A�9�*�LW�W� N�9�{�*�Zb���QCdCHK0�j�ݠnI_��M�JļR oh�Q ��sJ�-v㩾�S �$�X �1�N�I�RC�H_D$RN���^�LE��i��p�Zh8�ţMSW�FL/M�PSCRF�75�Ҽ ��3�" Ķ�6��`��ع�����0SV��Pp'������GRO�g�S_SA=AH�=��NO^`Ci�_d =��no�O�O�x�ʚ�`�p�B�u�ȐcDO�A��!�ں�*�tҀ:�Z1f�;�7����C ��Q�0Mmu� � �YL�snQ ��� ���"��<s�	�����nQ૰<N3M_Wl�����\p��(�o�MC��P���Q����rhpM.�pr� ��!ȅ�$�WM��ANGL�!�AM�6dK�=d@K�DdK��TT7�Nk@P��3�#�PXC OEc¼QZ��hp	nt� -���OM���� �ϣϵ����`� c�Z0��� L^a_�2� |a�J��i���c ���cJ��j�����jAB� ���{���  ��@{�P�1�PM�ON_QU�� �� 860QCOU���QTHxHO܆�B HYS�0ES�PBB UE- 3�f0O.�4�  c P�~^�RUN_TO���l�O��� P�@��INDE�#_PGRA���0��}2��NE_NO�ƋITf��o INFO��a"������P!OI� (*�SLEQ!�*��*�&S��l4�{ 460ENABy�>� PTION�3�p�r��^GCF�!� @60J�Q���R�d!���
�PEDIT�ԓ �� ��KAQ"�� �E(�NU'(A�UTY�%COPY�AQ�2,�qe�M�Nx< @+��PRUTm� C"N�OU�2�$G��$#RGAkDJ��u2X_��AIX����&���&W�(�P�(~��&9�� 
�N^�P_CYCy�H�/RGNSc�{�s��LGO£�NYQ__FREQSrW@��X1�4�L�@�2P0p�!�c@�"�CRE���MàIF�q�NA���%�4_Gf�S�TATU~�f��M'AIL��|CIq�=�LAST�1a*4EwLEMg� ��Q>rFEASIt;� ւΰ��B"�F�AF����I� ��O2�E� u�vBAB��PE� =�VA�FzQ�I��bTqU[��R��S~�FRMS_TRpC �Qc��C��Z�
��1�DX  *4ns؆�	MB? 2� `��� N�3V�R2WR*����p�R^W�wj�DOU�2^�N�,2PR`�h=�1GRID��oBARS!�TYu�Z�Op�� �|_�4!� �R�TO|��d� � ����POR�c~vb�SRV�0)"dfDI[�T�`;aNd�pXgD
�Xg4Vi��Xg6Vi%7Vi8:a�Fʒg��z $VALU��C0�3D��l�F05�� !pf���S1�1-ȆAN/��b��1R�]11ATOTcAL����=sPWE3�I�QStREGENQzfr��X�H�]5	�v( TR�CS�Qq_!S3��wfp�V�!��r��BE�3�PG0B��( sV_H�PDqA(��p�S_Ya����i6S��AR(�2�� �"IG_S!E�3�pb�5_� �t{C_�V$CMPl��DEp�G���I�šZ~�X��R�aEN�HANC.� �p Qr�2���I#NT9`cq�F����MASK�3�@OVRMP �PD�1-��W��c�U�l�_RF|�{�V�PSLGP�
g�9�j5��,��;pDpS���4��aU������TE����`���`k���Jx^�Y�y3IL_Mx40�s��p��TQ( �P��@����V.�C<��P_ �R�F�M]�V�1\�V1j�2y�2�j�3y�3j�4y�4 j���p۲������vܲIN�VIB8�P6�#��*�2&�22�U3&�32�4&�42���6�|�J�  �T $MC_FK `� �L>�J�х�1pMj�Iу��zS ���1���KEEP_HNADD���!鴓@�C��0 	��Q����
�O!��v ���p
�և
�REM!�	�Cq�RF�]��b�U�4e	�HPW�D  �SB�M���PCOLLAAB*�p��/q�2cIT/0��Q"NO1�FCALp⎵��� , �FLv�AO$SYN���M���Ck��RpUP_D�LY��zDEL�A9�Dq�2Y AD�(���QSKIPNO�� �`� O��cNT����c�P_�  ��׾ ��cp���q�� ���o`��|`�ډ`��@�`�ڣ`�ڰ`��9�!O�J2R0  �lX�@TR3H��1AH��� �H���7�RD�Cq��� � R"�R, 5��R�1��8E��5TRGE�_C��RFLG"���9W�5TSPC�1�UM_H��2TH�2N}Q�;� ?1� �;��Q>02 � D� ˈ<��@2_PC3W��S���1Y0L10_�Cw2��,��� � $\� U@�� V7�����0��VU\����� rd���C� +��7��DrZ Gs�RUVL1[��1h���10]�_�DS�������PK 11�� lڰ����q��AT?��$�Q [7�� ��K 5T����HOME� )��c2h�n�������3h����!3E *�c4h�hz�����&0`5h���	//-/?/Q'6h�b/t/�/�/�/�/
�7h��/�/??L'?9? ���!8h��\?n?�?�?�?�? �_S���� � �Aa{p�����+�_�Ed� aT=�nD4vnCIO�ҎII@`�O��_O�P�E�C.r���PO{WE	�� X@��f� �$$uCd�S����j@k��3�3� �@��SI��G�P0�QIRT�UAL�O
QAAV�M_WRK 2 �7U 0  �5Q�n_zXk_�] ��\	�P�]�_3�8P��_�_�Ve�\#m/o��Q5ojo|o�dHPBS��� 1Y� <Xo�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯�ݯ�bC$�AXLM��@���c  �d�IN����P+RE
�E�J�-�'_UP��[�7QHP?IOCNV_��k �	�Pr�US>��g�cIO)�V 1]U[P $E`��Q0ս9lҿ8P?�� � ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o�o�o�o�m�LAR�MRECOV �a��-���LMD/G ��ɰ��LM_IF  ���ை����z�v���%�6�, 
 6�_��r� ��������̍$w��� ׏��8�J�\�n�����NGTOL  �a� 	 A �  ��ț�PPI�NFO ={� <v����1��  I�3�a�"rP��� t��������ί���>�o����j�|��� ����Ŀֿ������0�B�PzPPLIC�ATION ?����+��HandlingTool ��� 
V9.30�P/04ǐM�
�88340�å�F90����202�ť�|�Ϭ�7DF3���M̎�NoneM��FRAM� �6��Z�_ACTI�VE�b  sï� � p�UTOMO�Dz�A���m�CH�GAPONL�� ���OUPLEDw 1ey� �������g�CURE�Q 1	e{  T*���	p��xw���#r�g���e�HN����{�HTTHK)Y��$r��\[�m� ���O�	�'�-�?�Q� c�u����������� ��#);M_q ������ %7I[m� ��/���/!/ 3/E/W/i/{/�/�/�/ ?�/�/�/??/?A? S?e?w?�?�?�?O�? �?�?OO+O=OOOaO sO�O�O�O_�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q��c���1�TO��|��p�DO_CLEA�N��n��NM  �� �B�T��f�x���%�DSPDgRYR��m�HI���@/�����,�>� P�b�t���������ίj�MAXa�ۄ�������Xۄ������p�PLUGG��܇�Ӯ��PRC��B�" ��ׯF�OK���^ȔSEGF��K�� �����.�����,�8>�v���LAPӟ� ��Ϥ϶��������π�"�4�F�X�j߯�T�OTAL�7���U�SENUӰ�� ����ߖ�1�RGDI_SPMMC����C����@@Ȓ��O�ѐ�����_STRING 1
�ۿ
�M��S�l�
A�_ITE;M1K�  nl�g� y������������ 	��-�?�Q�c�u����������I/O SIGNALE��Tryout� ModeL�I�np��Simul�atedP�Ou�tOVER�RА = 100�O�In cyc�lP�Prog� AborP�~��StatusN��	Heartbe�atJ�MH F�aul��Aler�	�������*<N`  ׃G�ׁY�c��� ��////A/S/e/ w/�/�/�/�/�/�/�/wWOR��G�-1� ?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO�cOuO�O�O�NPO E��@E;�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8oJo�BDEV�Nu`�O bo�o�o�o�o�o�o ,>Pbt�������PALT��E?�A�S� e�w���������я� ����+�=�O�a�s����GRI�G뽑 1������	��-�?� Q�c�u���������ϯ�����)�����R �a�՟;��������� ѿ�����+�=�O� a�sυϗϩϻ���O�PREG��y��� -�?�Q�c�u߇ߙ߫� ����������)�;��M�_�q����$AR�G_-0D ?	��������  	$���	[��]���������SBN_CONFIG���� ��CII�_SAVE  ���)���TCEL�LSETUP ���%  OME�_IO����%M�OV_Hn�����R�EPd�����UTO/BACKY���#�FRA:\��� ����)�'`rl ��&� 7�"� 24�/06{  09:_35:24������͓����� �+=Oas��������� �/1/C/U/g/y/�/ /�/�/�/�/�/	?�/ -???Q?c?u?�?�?p�ׁ  _��_\�ATBCKCTL.TM���?�?�?O\ O��INI�Y��-���MESSA�G9�GA)��RKODGE_Ds�<��zH�Ow`�O��PAUS��@ !��� ,,		�����O �G�O__#_%_7_q_ [_�__�_�_�_�_�_��_%o���D�@TSK  �M&,O���UPDT�@EGd��`�FXWZD_E�NBED��fSTApDE��e��XIS�?UNT 2��&��(�� 	 �0|} Z��0&? �<_ �/� K��Ppp�<�bp�p��8t}V��)q{|��t�� B=�|o���;9Յ�!{D�xp�Q��gMETc��2LfE� P qA�|hiA��A��B-��B�B�y��}�?yJ�?���?:�&@5�W�?U�s@����}SCRDCFG� 1�� ��z����� ԏ�����Q=��� H�Z�l�~�����	�Ɵ -����� �2�D���域���GR�`�`�O����0NA����	���_EDC@1�n�� 
 �%{-�0EDT-q�0���%�p��"���Q-���������x����  ����!2����*�R�bB����*�q���ϧ���3 bϮ�@Ͻϯd?����� =�O���sϏ�4.ߞ� {�����W���	�߱�?ߏ�5��j�G���΀#������}�6 ��6��Z�����Z�����I��7����� &��λ�&m����B��8^ҿ����	̀��9K�o��9*�w��	�S�`�;��CR�� ��B/T//�/���w//��РNO_D�EL����GE_U�NUSE���IG�ALLOW 1���2p(*S�YSTEM*�s�	$SERV_GqR�;B0�@REGK5�$m3�|B0NUMxp:�3�=PMU� >�uLAY�p�|�PMPAL|D@�5CYC10�.��>�0�>CULS�U�?�=�2�AM3L�OWDBOXORI�t5CUR_D@�=�PMCNV�6�D@10�>�@T4D�LI�`=O_9	*P�ROGRAJ4PG_MI�>�OP�AL�E_UPB�7_B>$FLUI_RESU�7p_z?��_�TMRY>h0�, �/�b�_�_o o2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v����������"LAL_OU�T 1;l���W?D_ABOR�0?�d�ITR_RTN�  ����g�N�ONSTOǠ��� 8CE_RIA3_I0��ۀ���ŀFCFG ���۔��_LI�MY22ګ �?  � 	i�J���<e�g��5��� 9��������
����u��PAQPG�P 1�@����Q�c�u�4�CK0�����C1��9��@����PC��CV��]*��d��l��s��P����C[٤m��vꭠ������� �C����-���?�ÂHE� ONFqI�Pq�G�G_P�@;1� �%� ������ǿٿ���ϾG�KPAUSaA1�ۃ �B�W� �Eσ�iϓϹϟ��� �������#�I�/�m���eߣ��M��NFoO 1"���� �7��ߖ��C� w�Bb?	��;ӛ8����,,MA�@��� ģ�C��Tp��1VC3�����"��3���3�E�ŀO��c�COLL/ECT_�"�[�����EN�@��y���nk�NDE��"��3�"1234?567890�� \1�� ��֕H&��)M�r�\,L�^���]+ ������������C  2�Vhz�� ����
c. @R�v����t����� ��>��IO !���q���u/�/�/�/C'[TR�2"'-(׀b^)
��.R�#R-x�*W� 9_MOR�$� �;�l5��l9 �?r?�?�?�?�;E2�*�%S=,W�?@�@�I�C׀K)DցC��R�&u�XOWAWBC�4  A&��׀x�׀A"@Cz  �B�@CG�B8��AC�  %��׀�ց:d�43 <#�
�E���I�OT�C=AI��'GM?�C��(S=���Qd=AT�_DEFPROG �;%�/m_APINUSE�V�ۅ��TKEY_TBL�  s�ہ���	
��� !"�#$%&'()*�+,-./�:;�<=>?@ABC�DPGHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����Ga���͓��������������������������������������������������?������!�P�LCK�\���P�PS�TAn��T_AUT/O_DO��NFs�IND���n��R_3T1wT2N�����5ŀTRLCPL�ETE���z_S�CREEN ~�kcscÂ�U��MMENU ;1)O� <�[_ #�q��,�a���>�d� ��t���ӏ����	��� ��Q�(�:���^�p� ������̟�ܟ�;� �$�q�H�Z������� ���Ưد%����4� m�D�V���z���ٿ�� ¿�!���
�W�.�@� ��d�vϜ��ϬϾ�� ����A��*�P߉�`� r߿ߖߨ�������� =��&�s�J�\��� ���������'�,�p_MANUAL��EqDB
12�v�iDBG_ERRLIPs*�{h! 0�������g�NUMLIM�s:QOE�@�DBPXWORK 1+�{��>P�bt��-DBTB_�q ,��kC3!�VD!DB_A�WAYo�h!GC�P OB=��A�_CAL���o�k�Y�p�uO@`�_�� 1-
�+@
-k-6[l��_M+pIS�`��@"@�ONTImM�w�OD���&
�U;MOTN�END�_:REC�ORD 13�{� ��[CG�O� f!T/[K��/�/�/�/ _(�/�/f/?�/??Q? c?�/?�??�?,?�? �?OO�?;O�?_O�? �O�O�O�O(O�OLO_ pO%_7_I_[_�O_�O �__�_�_�_�_l_!o �_,o�_io{o�o�oo �o2o�oVo/A �oeP^�
�� �R���=��a� s��������*�ߏN� ��'���ԏ]�̏�� ������ɟ۟v���n� #���G�Y�k�}����TOLERENC��B�0� L���g�CSS_CNS�TCY 24	�t���.����� �0�>�P�b�x����� ����ο����(��:�äDEVICEw 25ӫ � �ϟϱ������������/�AߟģHND�GD 6ӫ� C�zT�.!ơLS 27t�S������������/�U�ŢPARAM 8Gb��A�Ք�RBT 2]:8�<����CkA� �·�  � �A���.SB����A�B�  ����������.�����  ����A�A�C����c�u����C�A�D���k�pz�A�A��HA�c��A�	�?( uL^p���A��Bt/�D��C���_ 	 A�=��ABffA�#33AҊ��g�A�A�Cf���a��A�J��7B�]��B��B�ffBᴠ�3�3C$.@R� (����A��� �
/��//)/;/ �/_/q/�/�/�/�/�/ �/�/<??%?r?I?[? m??�?�?�?�?�?&O 8O�PObOMO�OqO�O �O�O�O�O_�OO L_#_5_�_Y_k_�_�_ �_�_ o�_�_6ooo loCoUogo�o�o�o�o �o�o �o	h�O �w�����
� �.�	__I'�1_� q��������ˏݏ� ��%�r�I�[���� ������ǟٟ&���� \�3�E�W����ȯ�� �ׯ�"��F�1�j� E�s�����m������� ѿ�0���f�=�O� a�sυϗ��ϻ���� ����'�9�Kߘ�o� ������[����(�� L�7�p��m��� ��������$����� l�C�U���y������� ���� ��	V-? �cu����
 ��@+dO�s ��������*/ //`/7/I/[/m// �/�/�/�/?�/�/? !?3?E?�?i?{?�?�? �?�?�?�?�?FO�jO UOgO�O�O�O�O�O�O __�'O9OO=_O_ �_s_�_�_�_�_�_�_ �_oPo'o9o�o]ooo �o�o�o�o�o�o: #5��O��� �� ��$��H�Fz��$DCSS_S�LAVE ;����w���`�_4D  �w���AR_MEN/U <w� >�؏@���� �2�^rǏ�\�n�\���SHOW� 2=w� � fr[q����Ə��� ��,�>�D�b�t��� ����ҟϯ��� �)�P�M�_�q����� ����˿ݿ���:� 7�I�[ς�|Ϧ��ϵ� ��������$�!�3�E� l�fߐύߟ߱����� �����/�V�P�z� w����������� ��@�:�d�a�s��� ��������\���*� H�N�K]o��� �����28� GYk}���� ��"�1/C/U/ g/y/�/��/�/�/� �//?-???Q?c?u? �/�?�?�?�/�??O O)O;OMO_O�?�O�O �O�?�O�?�O__%_ 7_I_pOm__�_�O�_ �O�_�_�_o!o3oZ_ Woio{o�_�o�_�o�o �o�oDo-Se �o��o�������.�=�O���CFoG >������q��dMC:�\��L%04d.'CSV\��pc����m���A ՃCH݀�z�v�w�#��q���:�J�8�7����JP�j�)�́�p+�n�RC_O�UT ?z����a�_C_F�SI ?�� |���� �@�;�M�_������� ��Я˯ݯ���%� 7�`�[�m�������� ǿ�����8�3�E� Wπ�{ύϟ������� �����/�X�S�e� wߠߛ߭߿������� �0�+�=�O�x�s�� ������������ '�P�K�]�o������� ����������(#5 Gpk}���� � �HCU g������� � //-/?/h/c/u/ �/�/�/�/�/�/�/? ?@?;?M?_?�?�?�? �?�?�?�?�?OO%O 7O`O[OmOO�O�O�O �O�O�O�O_8_3_E_ W_�_{_�_�_�_�_�_ �_ooo/oXoSoeo wo�o�o�o�o�o�o�o 0+=Oxs� �������� '�P�K�]�o������� ����ۏ���(�#�5� G�p�k�}�������ş ן �����H�C�U� g���������دӯ� �� ��-�?�h�c�u� ��������Ͽ���� �@�;�M�_ψσϕ� ������������%� 7�`�[�m�ߨߣߵ� ���������8�3�E� W��{��������� �����/�X�S�e� w��������������� 0+=Oxs� ����� 'PK]o��� �����(/#/5/ G/p/k/}/�/�/�/�/ �/ ?�/??H?C?U3��$DCS_C_�FSO ?�����1 P [?U?�?�? �?�?�?O
OO.OWO ROdOvO�O�O�O�O�O �O�O_/_*_<_N_w_ r_�_�_�_�_�_�_o oo&oOoJo\ono�o �o�o�o�o�o�o�o' "4Foj|�� �������G� B�T�f���������׏ ҏ�����,�>�g� b�t���������Ο�� ���?�:�L�^����������ϯʯܯg?C/_RPI~>�?� ;�d�_�
�}?.�p���X�ݿj>SL�@�� �9�b�]�oρϪϥ� �����������:�5� G�Y߂�}ߏߡ����� �������1�Z�U� g�y���������� ��	�2�-�?�Q�z�u� ������������
 )RM_q�� �����*% 7Irm��� ��/�ϛ�,�/ W/�/{/�/�/�/�/�/ �/???/?X?S?e? w?�?�?�?�?�?�?�? O0O+O=OOOxOsO�O �O�O�O�O�O___ '_P_K_]_o_�_�_�_ �_�_�_�_�_(o#o5o Gopoko}o�o�o�o�o �o �oHCU g��������� ����NOCO�DE @������PRE_?CHK B��3��A 3��< �7��������� 	 <�����?# ۏ%�7��[�m�G�Y� ������ٟ�ş�!� ���W�i�C�����y� ïկˏ������A� S�-�_���c�u���ѿ �������=��)� sυ�_ϩϻϕ����� ���'�9���E�o�I� [ߥ߷ߑ��������� #����Y�k�E��� {����������� C�U��=�����w��� ������	����?Q +u�a���� ��);_q g�Y��S��� �%/�/[/m/G/�/ �/}/�/�/�/�/?!? �/E?W?1?c?�?�� �?�?o?�?O�?�?AO SO-OwO�OcO�O�O�O �O�O_�O+_=__I_ s_M___�_�_�_�_�_ �?�_'o9oo]oooIo �o�oo�o�o�o�o #�oGY3E�� {�����o� C�U��y���e����� ������	��-�?�� K�u�O�a�������� �͟��)��1�_�q� �}�������ݯ�ɯ �%���1�[�5�G��� ��}�ǿٿ����� ��E�W�1�{ύ�G�u� ���ϯ������/�A� �-�w߉�c߭߿ߙ� ��������+�=��a� s�M���ϑ����� ���'��3�]�7�I� ������������� ����GY3}�i �������� C/y�e�� �����-/?// c/u/O/�/�/�/�/�/ �/�/?)?�?_?q? K?�?�?�?�?�?�?�? O%O�?IO[O5OO�O kO}O�O�O�O�O_�O 3_E_;?-_{_�_'_�_ �_�_�_�_�_�_/oAo oeowoQo�o�o�o�o �o�o�o+7a W_i_��C��� ��'��K�]�7�i� ��m��ɏۏ����� ��G�!�3�}���i� ��ş������1� C��g�y�S�e����� �����ѯ�-��� c�u�O�������Ͽ� ןɿ�)�ÿM�_�9� kϕ�oρ����Ϸ�� ����I�#�5�ߑ� kߵ��ߡ������� 3�E���Q�{�U�g�� ����������/�	� �e�w�Q��������� ������+Oa �I������ �K]7� �m�����/ �5/G/!/k/}/se/ �/�/_/�/�/�/?1? ??g?y?S?�?�?�? �?�?�?�?O-OOQO cO=OoO�O�/�/�O�O {O�O_�O_M___9_ �_�_o_�_�_�_�_o o�_7oIo#oUooYo ko�o�o�o�o�o�O�o 3Ei{U�� ������/�	� S�e�?�Q�������я ㏽����O�a� ������q���͟���� ���9�K�%�W��� [�m���ɯ�����ٯ �5�+�=�k�}���� ���������տ�1� �=�g�A�Sϝϯω� ���Ͽ�������Q��c����$DCS_SGN CS�����#M��27-JUN-�24 09:44� E�06��3�9������ /X�L��������������ДќM��Þ�j������{�VERSIO�N ��V�4.2.10�E�FLOGIC 1�DS��  	D���X�k��X�z�M�PROG_�ENB  ���b��Л�ULSE � ���M�_A�CCLIM��������WRS�TJNT����w�EMO���ѷ�L���INIT E�Z�O��OPT_�SL ?	S�1�
� 	R575��Ӆ�74��6��7R��5A��1��2���l���G�h�TO  �t���.H�V?�DKEX��d����FPATH A�ڇA\4���H�CP_CLNTI�D ?+�b� �l�����IAG_GRP 2JS�� ��a[�D�  �D�� D  �B�  B�@3ff��/B�@[���W�@�q���B�N�C�-Bz��Bp@�e`��mp�3m7 7890?123456�*��[��  Ao��mAj1Ad�A]�
AW�|�AP�AJ�-AC/A;��A4H���@��  A��A�A,3!_A�@@��;B4�� ��t����
�uƨAp�ffAj�yAe�K�A_�AYAS� MC��AF��A@ � O�+/=/O$O�c K�w(�@�X?8��@��y�/�/�/��/�/8�;d�2��5?@~ff@x�1'@q��@k�C�@d�D@]?��@Vv�6?H?�Z?l?~?8s�0l���@e@^���@W\)@O���@H�0?<@7K�@.V�?�?�?��?
O8S@M�00G<@A��@<�1@5��@/�l�@(Ĝ@!�0�\NO`OrO�O �Ox'g�L_K�;_�_�_ _g_�_�_�_�_o�_ �_�_YokoIo�o�o+o�oX�"� 2�17A��@J>��R
q?�33?Y��r���J7'Ŭz2q63p4�F>r���LJ@�p��Zr�
=@�O@�Q�jq��@G �Ah�@��@�T=� c<��]>�*�H>V>�3�>���J?<���<�p�q��x��� �?� ��C�  <(��U�� 4Vr�3a3��@
���A@��?R�oD��mR�x��� Q��t����Z�Џ��؏x�,��i?�7N��>�(�>�@Z�=����J��G�v�G�J�B�E������a��@ǐ@����@��@Q�?LT ���ŲI��P���&���' ��@�K����Ag�q�P�C�  C���CCuy�
���ʯ ?� ���	��Գ�4���X���v���*C�z�C�8�D��h�3��6C �F�ǿB���ֿ����E�T���� =�2�������=��^>��&$
�Iϗ�C�T_CONFIG� K3����eg��ST�BF_TTS��
@����"�������{��MAU���MS�W_CF��L � K �OCVIE�W	�MI�U�� 㯛߭߿��������� ���0�B�T�f�x�� ������������� ,�>�P�b�t������ ����������(: L^p���� �� �6HZ l~�����X�/��RCB�N��!��F/{/j/�/��/�/�/�/��SBL�_FAULT �O9*^�1GPMS�K��7��TDIAOG P��U�����qUD1�: 6789012345q2�q���%P�ϭ?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O �a6�I'��
�?_��TREC	PJ?\:
j4\_�7_[ �?�_�_�_�_�_�_o o(o:oLo^opo�o�o��o�o�O�O_ _�U�MP_OPTIO1N��>qTRB���:9;uPME��.�Y_TEMP  È�3B����p�A�pytUNI�'��ŏq6�YN_B�RK Qt�_�EDITOR q&qh��r_2PENT 1�R9)  ,&�COLOCA_�bpA_IRVIS�$r5� &MA�IN %�b�&�DROP_DEF}E�p_3 O ]���cv�2���v�1t��Ĉx�SEM|����Ɔ �BARR;A_�pNO ����&PEG-�E?STEIRA:����&PICKUUP��M�P�p 
����&SEGU�2�/����� &SUMIR ������ʂؓF��DA_?PRENSA�Ƀ1���8� A�ʂ���1_PLACqE0>�H�&
T�05�4�n���&ؓ/�����R���/�ǯy�b�4���٥�/����8�J��%EMGDI_STA�u�~��q�uNC_IN�FO 1SI��b�������Կⷮ�v��1TI� ��o#�Ϡ�0�d�o}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������Hu� �2� D�R�j�R�x���� ����������,�>� P�b�t����������� ��Z��#5Ga� k}������ �1CUgy ��������	/ /-/?/Yc/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?��?O%O7OQ/ GOmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�?O oo/o�_[Oeowo�o �o�o�o�o�o�o +=Oas��� ���_�_��'�9� So]�o���������ɏ ۏ����#�5�G�Y� k�}�������şן� ����1�K�U�g�y� ��������ӯ���	� �-�?�Q�c�u����� ����Ͽ����)� C�5�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ���� �����!�;�M�W�i� {������������ ��/�A�S�e�w��� ������������ +E�Oas��� ����'9 K]o����1 ����/#/=G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?��?�?	O O5/?OQOcOuO�O�O �O�O�O�O�O__)_ ;_M___q_�_�_�_�_ �?�_�_oo-O#oIo [omoo�o�o�o�o�o �o�o!3EWi {����_�_�� ��7oA�S�e�w��� ������я����� +�=�O�a�s������� ��ߟ���/�9� K�]�o���������ɯ ۯ����#�5�G�Y� k�}�������͟׿� ���'�1�C�U�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� ��ſ��������� ;�M�_�q����� ��������%�7�I� [�m�������߯��� �����)�3EWi {������� /ASew� ��������/! +/=/O/a/s/�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?/��? �?�?�?/#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�?�_�_�_�_O o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���_� ���	o�%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�����ß՟矝� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߩ��������� ���1�C�U�g�y� ������������	� �-�?�Q�c�u����� ������������) ;M_q���� ���%7I [m������ ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?S?e?w?� ��?�?�?�?�OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�?�?�_�_�_ �_�?�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �_�����_�	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q��y����� ˟�۟��%�7�I� [�m��������ǯٯ ����!�3�E�W�i���� �$ENETMODE 1U���  ��������»���RROR_PR_OG %��%������TABLE  ���Q�c��uσ��SEV_N�UM ��  �������_A�UTO_ENB � ̵��ݴ_NON�� V������_  *������%��������+���x(�:���FLTR����HIS�Ð�����_ALM 1W��� ����̍�+;���������0�r?�_����  �����²u꒰TCP_VER !���!��@�$EXTL�OG_REQv�9�����SIZ�����STK�����~��TOL  ��{Dz~��A ��_BWDU�*�Z�V��ǲ?�DID� X�Z�����[�STEPl�~�����OP_DO���F�ACTORY_T�UNv�d��DR_?GRP 1Y��`чd 	p�.° ��*u����RHB ��2 ���� �e9 ���bt�o ��������J5nYA����A'�q@9��u��
 J���ȸo��_�/�(/(B�  �F!A�  @�3�3R"�33-@UUTn*@P  /ȷ�>u.�>*���<��ǆ-E��� F@ �"�5�W�%�-J��NJ�k�I'PKH�u��IP�sF�!���-?�  �?�/9�<9��896C�'6<,5����-�YHv ��� �"�9d���A��FEATURE �Z�V�Ʊ�Handlin?gTool �5���Englis�h Dictio�nary�74D ;St�0ard�6�5�Analog I�/O�7�7gle �Shift Out�o Softwa�re Updat�e%Imatic ?Backup�9SA�ground E�dit�0�7Cam�era�0F�?Cn?rRndImXC�L�ommon ca?lib UI�C�F�nqA�@Monit�or�Ktr�0Re�liab@�8DH�CP�IZata ?Acquis�CY?iagnosOA�1�[ocument? Viewe�BW�ual Chec�k Safety��A�6hancedh�F�:�UsnPFr�@��7xt. DIO� �@fiRT�Wen]d�PErr�@LQR��]�Ws�Yr�0�P �E�:FCTN M�enu�Pv S8gT�P In'`fac<Ne�5GigE`nre�j@p Mask �Exc�Pg�WHT�^`Proxy S�voT�figh-S;pe�PSki�D�e�JP�PmmunicnN@ons�hurE`�'`_�1abconn�ect 2xnc=r``stru�2z�>peeQPJQU�4K�AREL Cmd7. L�`ua�hus�Run-Ti�PE�nvkx(`el +�R@sP@S/W�7L?icense�Sn\��PBook(Sy�stem)�:MA�CROs,�b/OOffse@�uH�P8@_�pMR�@�BP^�MechStop"�at.p6R�ui�RK�j�x�P�0P@)�od>@witch��>��EQ.���Optm8Џ>��`filn\=��gw�uulti-�T�`tC�9PCM 'funHwF�o3T�R�?�f�Regi�pr,�`I�rigPFV�����0Num Sel�b����P Adju��`���J�tat�u��
�iZ�5RDM� Robot�0s�cove�1F�ea�7��PFreq Awnly�gRem`���Qn�7F�R�Ser�vo�P���8SNPgX b�rNSN^`�ClifQɮBLi#br�3鯢0 q���굦o�ptE`ssag?��4�� -C��;��/I_mB�MIL�IBk�E�P Fi�rm6BU�PEcAcyck@sKTPTX_C�eln���F��1��V�orqu@i�mula�A�A�u��Pa�qU�j@�Ã�&�`ev.B�.@r�iP޿USB �port �@iP��PagP��R EV�NT�ϗ�nexcept�P��t��ſX�]VC�Ar�b�bf��V2PҦ�$����S�ܠSCصV�SGE�k�a�UI�;Web Pl!��ާ����`�TeQfZDT Appl�d�:�ƺ�� �GridV�plCay�R�WD4�R
��.�:n�EQ+��r-1?0iA/7L*��1Graphic��v�5dv�SDCSJ��ck�q�5larm Cause/���ed�8Ascii<�a��LoadnP�'Upl,�Ol�0�A�Gu�6N�`���yFyc@�r�����PV��3Jo��m� c�R��0�c���m�./����0�Q�2*u:eRAJ��P�ٶ4eqinL����8gNRT��9On�0e Hel�HJ�`o�I�alletiz`?�H�����_�tr�[ROS Eth�q��T@e�ׅ�!�n�%�;2D�tPkg&�Upg~�(2�DV-�3D T�ri-jQEAưD�ef.qEBa)pd�ei��� �bIm�πF�f��nsp�.q=�464MB �DRAMZ,#FR9O5/@ell�<�M#shf!r/�'c%�3@pLƖ,ty@s ˒xG��m��.[��  ��BU���Q�B�=mai�P߫�]Q����@q6wlu����^`��xR�?eL� Su�p������0�P�`cr��@�R���b䚮�p�r1uest�rt~QQ��ߋL!�4O��q$�K��l B�ui7�n��APL�COO�EVl%��CG�U�OCRG�O��D�R��O
TLS_��B�U/_��K�qN_d�T	A�OxVB�_�W�ܑZ���_TCB�_�V�_�W���WF+o�V�O�Wp._�W�ņoTEH�o`�f�O�gt�oTEj�BxVF�_w�_xVGo TwBTw~oxVH�xV�IA��v�xVLN�yUMz�bo�f_xVN�xVP���^xVR&xVS��܇ʏ���W��v���VGF:�L�P2_h�� h�V�h��_g�D��h�aFFoh��g�RD�n� TUT��01:��L�2V�L�TBGG���v�rain�U9I��
%HMI���Gpon��m�f��"�F�&KAR3EL9� �TPj���<6 SWIMESMTڢF0O�<5�
" a�X�j�������ͿĿ ֿ���'��0�]�T� fϓϊϜ��������� ��#��,�Y�P�bߏ� �ߘ��߼�������� �(�U�L�^���� �����������$� Q�H�Z���~������� ������ MD V�z����� �
I@R v������/ //E/</N/{/r/�/ �/�/�/�/�/??? A?8?J?w?n?�?�?�? �?�?�?O�?O=O4O FOsOjO|O�O�O�O�O �O_�O_9_0_B_o_ f_x_�_�_�_�_�_�_ �_o5o,o>okoboto �o�o�o�o�o�o�o 1(:g^p�� ����� �-�$� 6�c�Z�l��������� Ə����)� �2�_� V�h���������� ���%��.�[�R�d� �������������� !��*�W�N�`����� �������޿��� &�S�J�\ωπϒϤ� ����������"�O� F�X߅�|ߎߠ߲��� �������K�B�T� ��x���������� ���G�>�P�}�t� ������������ C:Lyp�� ����	 ? 6Hul~��� ��/�/;/2/D/ q/h/z/�/�/�/�/�/ ?�/
?7?.?@?m?d? v?�?�?�?�?�?�?�? O3O*O<OiO`OrO�O �O�O�O�O�O�O_/_ &_8_e_\_n_�_�_�_ �_�_�_�_�_+o"o4o aoXojo|o�o�o�o�o �o�o�o'0]T fx������ �#��,�Y�P�b�t� ������������� �(�U�L�^�p����� �����ܟ���$� Q�H�Z�l�~������� �د��� �M�D��V�h���  �H552}���2�1��R78��50ީ�J614��AT�UPͶ545͸6ީ�VCAM��CR�I�UIFͷ28n	�NRE��52��wR63��SCH���DOCV]�CSU���869ͷ0ضE�IOC9�4��R6=9��ESET����J7��R68��M�ASK��PRXY�!�7��OCO��3�帨���̸3�J6�˸53��H2�LC�H��OPLG�0^�MHCR��S{��MCS�0��55�ضMDSW���OP�MPR�M�@��0̶PCM �R0`���ض��@�51��51<�0�PRSv��69�FRD��FREQ��MCN���93̶SNBA�E�3�SHLB��M���M���2̶HTC��TMIL����T{PA��TPTX��#EL��Ѐ�8����J95,�TUTv�95�UEV��wUEC��UFR��VCC��O��VI�P�CSC,�CS�G8�r�I��WEBn�HTT�R6CȶN�CGIG��I�PGS)RC�D]G�H77��6ضwR85��R66��R7��R:�R53�0�680�2�q�JT��H�6<�6,�RJ�ԭ�0�4�6o64�\�5�NVD��R6��R84Tg�����8�90\���JM93�91� 7+Ǭ��,�D0oF�CsLI���CMS��� �STY��TOh�q���7�NN�ORS��J% ��j�OL(END��L���Sf(FVR��Vs3D���PBV,�wAPL��APV�wCCG�CCR|ֻCD��CDL@C�SBt�CSK��CT�CTBL9��U0�,(C��y0L8C��T�C �y0�'TC(7TC��CTE\��07cTEh��0��TFd8�F,(GL8GI�8H¸8I��E@�87�CTUM,(M�8M@8N�8�PHHPL8Rd8(T�Sd8W�I@VGF6�GP2��P2���@\�H{7VPD�HF ƻVPSGVPR�&VqT��YP��VTB7-Vs�IH��VI aH�'VK��VGene�����_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ �����/�A�S�e� w���������џ��� ��+�=�O�a�s��� ������ͯ߯��� '�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�?�  H5�5hT�1�1[U�3R7�8�<50�9J61�4�9ATU�T�45�45�<6�9VCA��D�3CRI,KUI�8T�528-JNREv�:52JR63�;�SCH�9DOCVr�JCU�4869�;�0�:EIO�TsE4�:R69JESE�T�;KJ7KR6�8�JMASK�9P�RXYML7�:OC�O\3�<�J)P�<3�|ZJ6�<53�JH�\LCH\ZOPL�G�;0�ZMHCR�]ZSkMCS�<0�,[55�:MDSW�}k�[OP�[MPR�Z�@�\0�:PCMLJR0�k)P�:)`�[[51K51|0J�PRS[69|ZF{RD<JFREQ�:�MCN�:93�:S�NBA}K�[SHLEB�zM�{�@ll2�:�HTC�:TMILܽ<�JTPA�JTPTX�EL�z)`�Kq8�;�0�JJ95\J�TUT�[95|ZU�EVZUEC\ZU�FR<JVCC��O�<jVIP,�CSCN\�CSGlJ�@I�9wWEB�:HTT�:�R6{L��CG{�I�G[�IPGS��R�C,�DG�[H77��<6�:R85�JR[66JR7[R|�R53{68|2��Z�@Jml,|6|6�\JR�\	P|4L�6��64��5�kNV�DZR6+kR84�<���IP,�8��90l���KJ9�\91��b̫7[KIP\JD0��F��CLI�lKC�MS�J9��:STYF,�TO�:�@�K7�L�NN|ZORS<jJة�MZZ|OLK�EN�D�:L�S��FV�R�JV3D,�KKP�BV\�APL�JA�PV�ZCCG�:C�CRjCD�CD�L̚CSB�JCS�K�jCTK�CTB��\���\�C�z��܍CL�TCLJ�l�T�C��TCZCTE�J��|�TE�J��<��TF��F\�G��G��l�Hl�I�z)�l�k�CTM\�M\�M���Nl�P,�P��R,��;�TS��W��̚�VGF��P2��P�2�z �VPD�FLJVP;�VP�R��VT�;� �JVkTB��V�KIH��VِM�<�VK,�V{�Gene�8�83 EWi{���� ���////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?a?s? �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qc u������� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�[�m������ ��ǟٟ����!�3� E�W�i�{�������ï կ�����/�A�S� e�w���������ѿ� ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3?�E?W?i?{?�7�0�STD�4LANG�4�9�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~��������� �2�D�V�R{BT�6OPTNm� �������Ǐُ��� �!�3�E�W�i�{���p����ß�5DPN�4 �����/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5߀G�Y�k�}ߏߡ߳�ted �4�8������ ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ������*�<�N�`��r���99���$�FEAT_ADD ?	��������  	 ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu������DEMO� Z��   ���}��'�� 0�]�T�f��������� ������#��,�Y� P�b������������ �����(�U�L�^� �����������ܯ� ��$�Q�H�Z���~� �������ؿ���  �M�D�Vσ�zόϦ� ���������
��I� @�R��v߈ߢ߬��� �������E�<�N� {�r���������� ���A�8�J�w�n� �������������� =4Fsj|� �����9 0Bofx��� ����/5/,/>/ k/b/t/�/�/�/�/�/ �/�/?1?(?:?g?^? p?�?�?�?�?�?�?�?  O-O$O6OcOZOlO�O �O�O�O�O�O�O�O)_  _2___V_h_�_�_�_ �_�_�_�_�_%oo.o [oRodo~o�o�o�o�o �o�o�o!*WN `z������ ���&�S�J�\�v� ���������ڏ�� �"�O�F�X�r�|��� ����ߟ֟���� K�B�T�n�x������� ۯү����G�>� P�j�t�������׿ο ����C�:�L�f� pϝϔϦ�������	�  ��?�6�H�b�lߙ� �ߢ����������� ;�2�D�^�h���� ���������
�7�.� @�Z�d����������� ������3*<V `������� �/&8R\� �������� +/"/4/N/X/�/|/�/ �/�/�/�/�/�/'?? 0?J?T?�?x?�?�?�? �?�?�?�?#OO,OFO PO}OtO�O�O�O�O�O �O�O__(_B_L_y_ p_�_�_�_�_�_�_�_ oo$o>oHouolo~o �o�o�o�o�o�o  :Dqhz�� �����
��6� @�m�d�v�������ُ Џ����2�<�i� `�r�������՟̟ޟ ���.�8�e�\�n� ������ѯȯگ��� �*�4�a�X�j����� ��ͿĿֿ����&� 0�]�T�fϓϊϜ��� ���������"�,�Y� P�bߏ߆ߘ��߼��� ������(�U�L�^� �������������  ��$�Q�H�Z���~� ��������������  MDV�z�� �����I @Rv���� ���//E/</N/ {/r/�/�/�/�/�/�/ �/
??A?8?J?w?n? �?�?�?�?�?�?�?O O=O4OFOsOjO|O�O �O�O�O�O�O__9_ 0_B_o_f_x_�_�_�_ �_�_�_�_o5o,o>o koboto�o�o�o�o�o �o�o1(:g^ p�������  �-�$�6�c�Z�l��� ����ϏƏ؏���)�  �2�_�V�h������� ˟ԟ���%��.� [�R�d�������ǯ�� Я���!��*�W�N� `�������ÿ��̿� ���&�S�J�\ω� �ϒϿ϶�������� �"�O�F�X߅�|ߎ� �߲���������� K�B�T��x���� ���������G�>��P�}�t���������  ������ "4FXj|�� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz���|��y  �x �q���&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t��������� ο����(�:�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������q�p�x���*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p���������������$FEAT_�DEMOIN  ��� ������INDEX����ILECO�MP [���B��8 �SETUP2 �\BL� � N w5_AP2BCK 1]B	?  �)���"�%����E � 	���5�Y�f ��B��x/ �1/C/�g/��/�/ ,/�/P/�/t/�/?�/ ??�/c?u??�?(?�? �?^?�?�?O)O�?MO �?qO O~O�O6O�OZO �O_�O%_�OI_[_�O __�_�_D_�_h_�_ �_
o3o�_Wo�_{o�o o�o@o�o�ovo�o /A�oe�o�� �N�r���=� �a�s����&���͏ \�񏀏���"�K�ڏ o�������4�ɟX�� ����#���G�Y��}�����0���ׯQ	� P� 2� *.cVRޯ(���*+��Q���W�{�e��PC�������FR6:D��ؾg�����T    �2����\� ��d�*.F��ϕ�	ó����o�ߓ�STM�9���ư%�"d��ψߓ�HU߻��Jש�f�x���GIF�A�L�-����ߑ���JPG����Lձ�0n�����JS�H�■��6���%
J�avaScriptt���CSe���K����v� %Cas�cading S�tyle She�ets��j�
AR�GNAME.DT'��O�\;��[��k|(k DISP*rUOп���� �
TPEI?NS.XML/��:\CcCus�tom Tool�bar��	PAS�SWORD����FRS:\�� �%Passwo�rd Config/c�Q/�J/�/�� �/:/�/�/p/?�/)? ;?�/_?�/�??$?�? H?�?l?�?O�?7O�? [OmO�?�O O�O�OVO �OzO_�O�OE_�Oi_ �Ob_�_._�_R_�_�_ �_o�_AoSo�_woo �o*o<o�o`o�o�o�o +�oO�os�� 8��n��'�� �]�����z���F� ۏj������5�ďY� k��������B�T�� x�����C�ҟg��� ����,���P������ ���?�ί�u���� (���Ͽ^�󿂿�)� ��M�ܿqσ�ϧ�6� ��Z�l�ߐ�%ߴ�� [����ߣߵ�D��� h�����3���W��� �ߍ���@����v� ���/�A���e���� ��*���N���r��� ��=��6s�& ��\��'� K�o��4� X���#/�G/Y/ �}//�/�/B/�/f/ �/�/�/1?�/U?�/N? �??�?>?�?�?t?	O �?-O?O�?cO�?�OO�(O�O�F�$FIL�E_DGBCK �1]���@��� < ��)
SUMMA�RY.DG�OsL�MD:�O;_@�Diag Sum�mary<_IJ
C?ONSLOG1__�&Q_�_NQCon�sole log��_HK	TPACC�N�_o%o?oJU�TP Accou�ntin�_IJF�R6:IPKDM�P.ZIPsowH
��o�oKU[`Exception�oyk'P�MEMCHECK�5o�_*_K�QMe�mory Dat�aL�FUl�)6qRIPE�_$6��Zs%�q Packet L�_��DL�$�	r�qS�TAT���S�� %�rSta�tusT��	FTAP���:���Vw�Q�mment TB�D؏� >I)ETHERNE�ఏ
q�[�NQEt�hern�p�Pfi�gura�oODDCSVRF̏��ď�ݟd��� verify all���{D�.���DIF�F՟��͟b��s��d�iffd��
q��CHG01Y�@�R�篰f�z���-?��2 ݯį֯k�v������3a�H�Z�� ���ϥ�VTRNDIAG.LS��̿޿s�^q3� O�pe���q SQno�stic�w�ɿ)VDEV7�D�ATt�Q�c�u�g��Vis��Devisce�Ϫ�IMG7 �o����y��s�I�magߨ�UP���ES��T�FR�S:\�� �OQU�pdates L�ist �IJg�FLEXEVENQ��X�j߃�f�F� UIF Ev���B�,�s�)
PS�RBWLD.CM���sL������PP�S_ROBOWE�L��GLo�GRAPHICS4Dy��b�t��%4D� Graphic?s Fileu��A�Oɿ�rGIG����u�
YvGi�gE�ة�BN�?� )��HADO�W�����\sS�hadow Ch�ang���v2b~QRCMERR��n�\s� CFG Error��tail� MA���CMSGLIB��"^�o� ��T�)�ZD����/nXwZD6 ad�zHPNOTI����
/�/ZuNot�ific��H/��AGUO�/yO?�O'? P?OOt??�?�?9?�? ]?�?O�?(O�?LO^O �?�OO�O5O�O�OkO  _�O$_6_�OZ_�O~_ �__�_C_�_�_y_o �_2o�_?oho�_�oo �o�oQo�ouo
�o @�odv�)� M�����<�N� �r������7�̏[� �����&���J�ُW� �����3�ȟڟi��� ��"�4�ßX��|��� ���A�֯e����� 0���T�f�������� ��O��s��ϩ�>� Ϳb��oϘ�'ϼ�K� ���ρ�ߥ�:�L��� p��ϔߦ�5���Y��� }���$��H���l�~� ��1�����g����  �2���V���z�	��� ��?���c���
��. ��Rd����� M�q�<� `���%�I� �/�8/J/�n/ ��/!/�/�/W/�/{/ ?"?�/F?�/j?|??�?/?�?�?�$FI�LE_FRSPRT  ���0����8�MDONLY 1�]�5�0 
 ��)MD:_V�DAEXTP.Z�ZZ�?�?_OnK�6%NO Ba�ck file <9O�4S�6Pe?�O OO�O�?�O__?>_�O b_t__�_'_�_�_]_ �_�_o(o�_Lo�_po �_}o�o5o�oYo�o  �o$�oHZ�o~ ��C�g��	� 2��V��z������ ?�ԏ�u�
���.�@�~�4VISBCKH|A&C*.VDA�|����FR:\Z��ION\DATA�\v����Vision VD�B ��ŏ���'�5��Y� �j������B�ׯ� x����1���үg��� ����X���P��t��� Ϫ�?�οc�u�ϙ� (Ͻ�L�^��ς��)� ��M���q� ߂ߧ�6� ��Z�����%��I��������:LUI_�CONFIG �^�5m��� '$ h�F{�5������)�;�I���|xq�s����������� a��� $6��G l~���K�� � 2�Vhz ���G���
/ /./�R/d/v/�/�/ �/C/�/�/�/??*? �/N?`?r?�?�?�??? �?�?�?OO&O�?JO \OnO�O�O)O�O�O�O �O�O_�O4_F_X_j_ |_�_%_�_�_�_�_�_ o�_0oBoTofoxo�o !o�o�o�o�o�o�o ,>Pbt�� ������(�:� L�^�p��������ʏ ܏���$�6�H�Z� l��������Ɵ؟� ��� �2�D�V�h��� ������¯ԯ�}�
� �.�@�R�d������� ����п�y���*� <�N�`����ϖϨϺ� ����u���&�8�J� ��[߀ߒߤ߶���_� �����"�4�F���j� |������[����� ��0�B���f�x��� ������W����� ,>��bt��� �O��(:>�  xFS��$FLUI_D�ATA _�������uRESULT� 2`�� ��T�/wi�zard/gui�ded/step�s/Expert b��//+/=/O/�a/s/�/�/�*�C�ontinue �with G�ance�/�/�/?? (?:?L?^?p?�?�?�?� T-U��90 �� �?��6�9��ps�?0O BOTOfOxO�O�O�O�O �O�O�O� �_/_A_ S_e_w_�_�_�_�_�_��_�_n�?�?�?�<Frip�Oo�o �o�o�o�o�o�o! 3E_i{��� ������/�A�@S�o$on�HoAO��TimeUS/DST[������ +�=�O�a�s������'?Enabl�/˟ ݟ���%�7�I�[�Pm������T�?`{�ݯ����Æ24Ώ 3�E�W�i�{������� ÿտ翦����/�A� S�e�wωϛϭϿ��� ���ϴ�Ưد� G�~�Region�� �ߙ߽߫����������)�;�+Americasou��� �����������)�;��?�y�#߅�G�|Y��ditorL� ������#5GY�k}��+ Tou�ch Panel� �� (reco/mmen�)�� �*<N`r��U��e�w����|����accesd� ./@/R/d/v/�/�/�/�/�/�/Q|Con�nect to Network�/ (?:?L?^?p?�?�?�?��?�?�?�?Y���������!/��I�ntroduct s߆O�O�O�O�O�O�O __(_:_U^_p_�_ �_�_�_�_�_�_ oo$o6oHo e�Oeo ?O�X_�o�o�o�o '9K]o�� R_������#��5�G�Y�k�}�����h`�ooj}oߏ�o� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ쯫���Ϗ1�� X�j�|�������Ŀֿ �����0��A�f� xϊϜϮ��������� ��,�>���_�!��� E��߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~���O߱�s� ������ 2DV hz������ ��
.@Rdv ��������/ ��'/���`/r/�/�/ �/�/�/�/�/??&? 8?�\?n?�?�?�?�? �?�?�?�?O"O4O� UO/yO�OO?�O�O�O �O�O__0_B_T_f_ x_�_I?�_�_�_�_�_ oo,o>oPoboto�o EO�OiO�o�o�O (:L^p��� ����_ ��$�6� H�Z�l�~�������Ə ؏�o�o�o�/��oV� h�z�������ԟ� ��
��.��R�d�v� ��������Я���� �*��������C� ����̿޿���&� 8�J�\�nπ�?��϶� ���������"�4�F� X�j�|ߎ�M�_�q��� ������0�B�T�f� x����������� ��,�>�P�b�t��� �����������߱��� %��L^p��� ���� $�� 5Zl~���� ���/ /2/��S/ w/9�/�/�/�/�/ �/
??.?@?R?d?v? �?�/�?�?�?�?�?O O*O<ONO`OrO�OC/ �Og/�O�/�O__&_ 8_J_\_n_�_�_�_�_ �_�_�?�_o"o4oFo Xojo|o�o�o�o�o�o �O�o�O�O�oTf x������� ��,��_P�b�t��� ������Ώ����� (��oI�m��C��� ��ʟܟ� ��$�6� H�Z�l�~�=�����Ư د���� �2�D�V� h�z�9���]���ѿ�� ��
��.�@�R�d�v� �ϚϬϾ��Ϗ���� �*�<�N�`�r߄ߖ� �ߺ��ߋ�տ����#� �J�\�n����� ���������"���F� X�j�|����������� ���������� u7������ ,>Pbt3� ������// (/:/L/^/p/�/AS e�/��/ ??$?6? H?Z?l?~?�?�?�?�? ��?�?O O2ODOVO hOzO�O�O�O�O�O�/ �/�/_�/@_R_d_v_ �_�_�_�_�_�_�_o o�?)oNo`oro�o�o �o�o�o�o�o& �OG	_k-_��� �����"�4�F� X�j�|������ď֏ �����0�B�T�f� x�7��[����� ��,�>�P�b�t��� ������ί����� (�:�L�^�p������� ��ʿ��뿭��џӿ H�Z�l�~ϐϢϴ��� ������� �߯D�V� h�zߌߞ߰������� ��
��ۿ=���a�s� 7ߚ���������� �*�<�N�`�r�1ߖ� ����������& 8J\n-�w�Q� �����"4F Xj|������ ��//0/B/T/f/ x/�/�/�/�/�� �/?�>?P?b?t?�? �?�?�?�?�?�?OO �:OLO^OpO�O�O�O �O�O�O�O __�/�/ �/?i_+?�_�_�_�_ �_�_�_o o2oDoVo ho'O�o�o�o�o�o�o �o
.@Rdv 5_G_Y_�}_��� �*�<�N�`�r����� ����yoޏ����&� 8�J�\�n��������� ȟ�����4�F� X�j�|�������į֯ ����ˏ�B�T�f� x���������ҿ��� ��ٟ;���_�!��� �Ϫϼ��������� (�:�L�^�p߁ϔߦ� �������� ��$�6� H�Z�l�+ύ�Oϱ�s� ������� �2�D�V� h�z������������� ��
.@Rdv ����}���� ���<N`r�� �����//�� 8/J/\/n/�/�/�/�/ �/�/�/�/?�1?� U?g?+/�?�?�?�?�? �?�?OO0OBOTOfO %/�O�O�O�O�O�O�O __,_>_P_b_!?k? E?�_�_{?�_�_oo (o:oLo^opo�o�o�o �owO�o�o $6 HZl~���s_ �_�_���_2�D�V� h�z�������ԏ� ��
��o.�@�R�d�v� ��������П���� ����]������ ����̯ޯ���&� 8�J�\���������� ȿڿ����"�4�F� X�j�)�;�M���q��� ������0�B�T�f� xߊߜ߮�m������� ��,�>�P�b�t�� ����{ύϟ���� (�:�L�^�p������� �������� ��6 HZl~���� �����/��S �z������ �
//./@/R/d/u �/�/�/�/�/�/�/? ?*?<?N?`?�?C �?g�?�?�?OO&O 8OJO\OnO�O�O�O�O u/�O�O�O_"_4_F_ X_j_|_�_�_�_q?�_ �?�_�?�_0oBoTofo xo�o�o�o�o�o�o�o �O,>Pbt� ��������_ %��_I�[������� ��ʏ܏� ��$�6� H�Z�~�������Ɵ ؟���� �2�D�V� �_�9�����o�ԯ� ��
��.�@�R�d�v� ������k�п���� �*�<�N�`�rτϖ� ��g�����������&� 8�J�\�n߀ߒߤ߶� �������߽�"�4�F� X�j�|�������� �����������Q�� x��������������� ,>P�t� ������ (:L^�/�A�� e���� //$/6/ H/Z/l/~/�/�/a�/ �/�/�/? ?2?D?V? h?z?�?�?�?o�� �?�O.O@OROdOvO �O�O�O�O�O�O�O�/ _*_<_N_`_r_�_�_ �_�_�_�_�_o�?#o �?Go	Ono�o�o�o�o �o�o�o�o"4F Xio|����� ����0�B�T�o u�7o��[o��ҏ��� ��,�>�P�b�t��� ����iΟ����� (�:�L�^�p������� e�ǯ��믭���$�6� H�Z�l�~�������ƿ ؿ����� �2�D�V� h�zόϞϰ������� �Ϸ��ۯ=�O��v� �ߚ߬߾�������� �*�<�N��r��� �����������&� 8�J�	�S�-�w���c� ��������"4F Xj|��_��� ��0BTf x��[������ ��/,/>/P/b/t/�/ �/�/�/�/�/�/�? (?:?L?^?p?�?�?�? �?�?�?�?���� EO/lO~O�O�O�O�O �O�O�O_ _2_D_? h_z_�_�_�_�_�_�_ �_
oo.o@oRoO#O 5O�oYO�o�o�o�o *<N`r�� U_������&� 8�J�\�n�������co uo�o鏫o�"�4�F� X�j�|�������ğ֟ 蟧���0�B�T�f� x���������ү��� ���ُ;���b�t��� ������ο���� (�:�L�]�pςϔϦ� �������� ��$�6� H��i�+���O����� ������� �2�D�V� h�z���]������� ��
��.�@�R�d�v� ����Y߻�}����ߣ� *<N`r�� �������& 8J\n���� �����/��1/C/ j/|/�/�/�/�/�/ �/�/??0?B?f? x?�?�?�?�?�?�?�? OO,O>O�G/!/kO �OW/�O�O�O�O__ (_:_L_^_p_�_�_S? �_�_�_�_ oo$o6o HoZolo~o�oOO�OsO �o�o�O 2DV hz������ �_
��.�@�R�d�v� ��������Џ⏡o�o �o�o9��o`�r����� ����̟ޟ���&� 8��\�n��������� ȯگ����"�4�F� ��)���M���Ŀֿ �����0�B�T�f� xϊ�I����������� ��,�>�P�b�t߆� ��W�i�{��ߟ��� (�:�L�^�p���� ����������$�6� H�Z�l�~��������� ��������/��V hz������ �
.@Qdv �������/ /*/</��]/�/C �/�/�/�/�/??&? 8?J?\?n?�?�?Q�? �?�?�?�?O"O4OFO XOjO|O�OM/�Oq/�O �/�O__0_B_T_f_ x_�_�_�_�_�_�_�? oo,o>oPoboto�o �o�o�o�o�o�O�O %7�_^p��� ���� ��$�6� �_Z�l�~�������Ə ؏���� �2��o; _���K��ԟ� ��
��.�@�R�d�v� ��G�����Я���� �*�<�N�`�r���C� ��g���ۿ����&� 8�J�\�nπϒϤ϶� ���ϙ����"�4�F� X�j�|ߎߠ߲����� ������˿-��T�f� x������������ ��,���P�b�t��� ������������ (:����A� ���� $6 HZl~=���� ���/ /2/D/V/ h/z/�/K]o�/� �/
??.?@?R?d?v? �?�?�?�?�?��?O O*O<ONO`OrO�O�O �O�O�O�O�/�O�/#_ �/J_\_n_�_�_�_�_ �_�_�_�_o"o4oE_ Xojo|o�o�o�o�o�o �o�o0�OQ_ u7_������ ��,�>�P�b�t��� Eo����Ώ����� (�:�L�^�p���A�� eǟ��� ��$�6� H�Z�l�~�������Ư د����� �2�D�V� h�z�������¿Կ�� �����+��R�d�v� �ϚϬϾ�������� �*��N�`�r߄ߖ� �ߺ���������&� �/�	�S�}�?Ϥ�� ���������"�4�F� X�j�|�;ߠ������� ����0BTf x7��[����� ,>Pbt� �������// (/:/L/^/p/�/�/�/ �/�/����!?� H?Z?l?~?�?�?�?�? �?�?�?O O�DOVO hOzO�O�O�O�O�O�O �O
__._�/�/?s_ 5?�_�_�_�_�_�_o o*o<oNo`oro1O�o �o�o�o�o�o& 8J\n�?_Q_c_ ��_���"�4�F� X�j�|�������ď�o Տ����0�B�T�f� x���������ҟ�� ���>�P�b�t��� ������ί���� (�9�L�^�p������� ��ʿܿ� ��$�� E��i�+��Ϣϴ��� ������� �2�D�V� h�z�9��߰������� ��
��.�@�R�d�v� 5ϗ�Yϻ�}����� �*�<�N�`�r����� ����������& 8J\n���� ��������F Xj|����� ��//��B/T/f/ x/�/�/�/�/�/�/�/ ??�#�G?q?3 �?�?�?�?�?�?OO (O:OLO^OpO//�O�O �O�O�O�O __$_6_ H_Z_l_+?u?O?�_�_ �?�_�_o o2oDoVo hozo�o�o�o�o�O�o �o
.@Rdv ����}_�_�_�_ ��_<�N�`�r����� ����̏ޏ�����o 8�J�\�n��������� ȟڟ����"��� �g�)�������į֯ �����0�B�T�f� %���������ҿ��� ��,�>�P�b�t�3� E�W���{������� (�:�L�^�p߂ߔߦ� ��w����� ��$�6� H�Z�l�~������ ��������2�D�V� h�z������������� ��
-�@Rdv ������� ��9��]��� �����//&/ 8/J/\/n/-�/�/�/ �/�/�/�/?"?4?F? X?j?)�?M�?qs? �?�?OO0OBOTOfO xO�O�O�O�O/�O�O __,_>_P_b_t_�_ �_�_�_{?�_�?oo �O:oLo^opo�o�o�o �o�o�o�o �O6 HZl~���� �����_o�_;� e�'o������ԏ� ��
��.�@�R�d�# ��������П���� �*�<�N�`��i�C� ����y�ޯ���&� 8�J�\�n��������� u�ڿ����"�4�F� X�j�|ώϠϲ�q��� ����	�˯0�B�T�f� xߊߜ߮��������� �ǿ,�>�P�b�t�� ������������ ������[�߂����� �������� $6 HZ�~���� ��� 2DV h'�9�K��o��� �
//./@/R/d/v/ �/�/�/k�/�/�/? ?*?<?N?`?r?�?�? �?�?y�?��?�&O 8OJO\OnO�O�O�O�O �O�O�O�O_!O4_F_ X_j_|_�_�_�_�_�_ �_�_o�?-o�?QoO xo�o�o�o�o�o�o�o ,>Pb!_� �������� (�:�L�^�o�Ao�� eog�܏� ��$�6� H�Z�l�~�������s ؟���� �2�D�V� h�z�������o�ѯ�� ���˟.�@�R�d�v� ��������п���� ş*�<�N�`�rτϖ� �Ϻ����������� �/�Y���ߒߤ߶� ���������"�4�F� X��|�������� ������0�B�T�� ]�7߁���m������� ,>Pbt� ��i���� (:L^p��� e�w��������$/6/ H/Z/l/~/�/�/�/�/ �/�/�/� ?2?D?V? h?z?�?�?�?�?�?�? �?
O���OO/vO �O�O�O�O�O�O�O_ _*_<_N_?r_�_�_ �_�_�_�_�_oo&o 8oJo\oO-O?O�ocO �o�o�o�o"4F Xj|��__�� ����0�B�T�f� x�������moϏ�o� �o�,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ���!�� E��l�~�������ƿ ؿ���� �2�D�V� �zόϞϰ������� ��
��.�@�R��s� 5���Y�[�������� �*�<�N�`�r��� ��g���������&� 8�J�\�n�������c� ����������"4F Xj|����� ����0BTf x������� ������#/M/t/�/ �/�/�/�/�/�/?? (?:?L?p?�?�?�? �?�?�?�? OO$O6O HO/Q/+/uO�Oa/�O �O�O�O_ _2_D_V_ h_z_�_�_]?�_�_�_ �_
oo.o@oRodovo �o�oYOkO}O�O�o�O *<N`r�� ������_�&� 8�J�\�n��������� ȏڏ����o�o�oC� j�|�������ğ֟ �����0�B��f� x���������ү��� ��,�>�P��!�3�������$FMR2_GRP 1a���� �C4  B�[�	 [�߿�ܰ�E�� F@ �5W�S�ܰJ���NJk�I�'PKHu��IP�sF!��͏?�  W�S�ܰ9��<9�8�96C'6<,5����A�  �Ϲ�BH�ٳB�հ����@ӻ33�33S��۴��ܰ@UUT�'�@��8��W�>u�.�>*��<�����=[�B=����=|	<��K�<�q�=��mo���8��x	7H<8��^6�Hc7��x?�����������"��F�X���_C�FG b»T �Q����X�N�O º
F�0�� ��W�RM_�CHKTYP  ���[�ʰ̰����R{OM�_MIN�[���9����X���SSBh�c��? ݶf��[�]����^�TP__DEF_O�[��ʳ��IRCOM����$GENO�VRD_DO.��d���THR.� dzd��_ENB��{ ��RAVC��udO�Z� ����Fs  G!� �GɃ�I�C��I(i J���+���%����ʷ �QOU��j�¼������<6�i�C�;]��[�C�  D0�+��@���B����.��R SMT��k_	ΰ\����$HOSTC�h�1l¹[��\d�۰ MC[����/Z�  2�7.0� 1�/  e�/??'?9?G: �/j?|?�?�?�,Z?T3�	anonymouy �?�?	OO-O?N�/ڰRHRK�/�?�O �/�O�O�O�O_V?3_ E_W_i_�O&_�?�_�_ �_�_�_@O�_dOvOSo �_�Ojo�o�o�o�o_ �o+=`o�_�_ �����o&o8o JoL9��o]�o����� ���oɏۏ����4� j+�Y�k�}������ ��� ��T�1�C� U�g�����������ӯ ��x�>��-�?�Q�c� ����Ο���Ͽ�� ��)�;ς�_�qσ� �ϧ�ʿ ������ %�7�~�����߶ϣ� ����������Ϻ�3� E�W�i�ߍ��ϱ��� ������@�R�d�v�x� J��߉���������� ��+=`�������:$h!E�NT 1m sP!V  7 ?.c&�J �n���/�)/ �M//q/4/�/X/j/ �/�/�/�/?�/7?�/ ?m?0?�?T?�?x?�? �?�?O�?3O�?WOO {O>O�ObO�O�O�O�O �O_�OA__e_(_:_��_^_�_�_�_�ZQUICC0�_�_�_?od1@oo.o�od�2�olo~o�o!ROUTER�o�o�o�/!PCJOG�0!192�.168.0.1�0	o�SCAMPRYT�\!pu1yp��vRT�o���� !Softw�are Oper�ator Pan�el�mn��NA�ME !�
!�ROBO�v�S_�CFG 1l�	� �Au�to-start{ed'�FTP2��I�K2��V�h� z�������ԟ��� �	���@�R�d�v��� 	�������:��� )�;�M�_�&������� ��˿�p���%�7� I�[��"�4�F�ڿ�� ������!�3���W� i�{ߍߟ���D����� ����/�vψϚ�w� �ߛ��Ͽ�������� �+�=�O�a������ ����������8�J�\� n�p�]����� �����#5X �k}���� 0/D1/xU/g/ y/�/RH/�/�/�/�/ /?�/??Q?c?u?�? ���/?�?:/O )O;OMO_O&?�O�O�O �O�O�?pO__%_7_ I_[_�?�?�?t_�O�_ O�_�_o!o3o�OWo io{o�o�_�oDo�o�o��o����_ER�R n��-=vP�DUSIZ  j�`^�P�Tt>mu?WRD ?΅�Q��  guest�f�������~�SCDMNGRP 2o΅wWp��Q�`���fKL� 	�P01.05 8~�Q   �|���  ;|���  z[ ����w���*����Ť�x�������[ݏȏ���ʑPԠ������)/����D�r��ꉫ؊p"�Pl�P���Dx��dx�*���|��%�_GROU7�UpLyN��	/�\o���QUP��U�Tu� �TYà�L}?pTTP_A�UTH 1qL{� <!iPen'dan����o֢�!KAREL:q*������KC���ɯۯ��VISI?ON SET�9� ���P�>�h��f��� �������ҿ�����X�CTRL �rL}O�uſa
��g�FFF9E3�-ϝTFRS:D�EFAULT���FANUC W�eb Server�ʅ�t�X���t@̀��1�C�U�g�;tW�R_CONFIGw s;� ���=qIDL_CPU�_PC���aB�ܠP�� BH��MI�N�܅q��GNR_�IOFq{r�`Rx��N�PT_SIM_D�O��STAL�_SCRN� ��.�INTPMOD�NTOLQ����R�TY0����-�\�E�NBQ�-���OL_NK 1tL{�p ������)�;�M���MASTE�%����SLAVE u�L|�RAMCAC�HEk�c�O^�O_�CFG������UO�C�����CMT_O�P���PzYCL�������_ASG s1v;��q
 O� r������� &8J\W�EWNUMzsPy
���IP����RTRY_CN��M�=�zs����Tu �������w���p/�p��P_�MEMBERS �2x;�l� $��X"��?�Q'W/i)���RCA_ACC �2y�  Xۿfn ��$�b6���"  0�` ���&�#�#�/�!���,��$BUF001 �2z�= c5�u� u0cG:4V�:4h:4x:4�:4��:4�:4�:4�:4�J:4�:3d=0�2�4U!�41�4C�4T�4eg�4w�4a4d��4U��4��4ђ4�4��:3e
D
D+�
D;
DN
Da
Dr�
D�
D�
D�
D��
D�4e�
D�:3fUzDzD&zD7zD�JzD[zDnzD�a   a bl:3�b|�D��D��D���D��D�4b��D�*:4:4:4%:392$?63:1@1ERI0ER Q0ERY0ERa0ERi0ER q0ERy0ER�0ER�0ER �0:1�1�R�0�R�0�R �0�R�0�R�0�R�0�R �0�RjT�1�R�0�R�0 �R�0�R@�R	@:1A b@b!@b)@b1@ b9@bA@bI@bQ@ bY@ba@b�TpAb y@:1�A�b�@�b�@�b �@�b�@�b�@�b�@�b�@(I��A:1�A �b�@�b�@�b�@�b�@ �bd�A�bPER	PER PERP:193-_65 GSNrI2WSNrY2gSNr i2wSNry2�SNr�2�S ���t�2�S���2�S�� �2�S���2�S���2�S ���2�S��Bc��C c�!B/c�1B?c� ABOc�QB_c�aBoc �qBc���C�c���B �c���B�c���B�c�� �C�c΂�B�c΂�B�c ΂��CsNr	RsNrXR'v��2{�4r�}ŋ���<����o��o��2�HIS!2}�� ܷ! 2�024-06-2�7����П��� � 8�;  X
�` 
�� m�)�;�M�_�o�/X�g��6�������Ư��o��o��g�#��"�4�F�}��j���5��~�������� 7 �h
�j�������.y��cN��1O�p��]�oρ� � 9 �cP��������\ ���mv��0��`5�G�Y�د�Z�M g9 ٰ��mvR��;�С߳�����`� ��!-��,�>�P�b� t���������� ��(�:�L�^�p��� ����,P����'�����Hoں�c���d�9� o�d_q� q��������q�I �I>��I6HZ lZ�l����!3:��b>ٰ9�9 �/1/C/1�C�L/�/��/�/
�� a >��	/�/ ??$?��Z?l?~?l�& S @6��;��c����o�c�?�?�?�? ����OCOUOgOyO�O �O�O�O�O
OO.O_ -_?_Q_c_u_�_�_�_ ����5p����L?o$o6oo��Td�VbF  Vbro�o�o�o��o �oKo]k��no[ m�����l�3t���ٰ2r �J?�Q�c�Q/c/� ����Ϗt��B��B�&�N����*�<� *?<?��������q�4sDp����֒���� ��
���O�Ow�d�v� ��������Я���� =�O�<�N�`�r�����ਿ��̿޿��I_C�FG 2~�[ �H
Cycle� Time�B�usy�Idl���min��S�Up���Read(�D�owG�Cϟ���Count�	ONum �������p�����PROmG���U�P��)/softp�art/genl�ink?curr�ent=menu�page,1133,1�C�U�g�y��Tä�SDT_IS�OLC  �Y�� ���J23_�DSP_ENB � ��T���INC� ���p���A �  ?�  =�?��<#�
���:�o �2�D�p�/�l���OB��C���O��ֆ�G_GROUP 1���;<*��(���t�?����p�Q'�L�^�p�/�����������\�~�G�_IN_AUTO|����POSRE�����KANJI_M�ASK0��DRELMON ��[��p�y������P��f�Ã�����p�-��KCL;_L NUM��G�$KEYLOGG'INGD�P��!�����LANGUAG�E �U���DEFAUL�T ��QLG��Y���S��p�x���ܐ8T�H  �p�'0��p��!֒�K�p�;��
*!(?UT1:\ J/ L/Y/k/}/�/�/@�/�/�/�/�/$>(��H?�VLN_DISP ���P�&�$��^4OCTOL�D�z����
�1GBO_OK ��d4V�11�0˕%O !O3OEOWOiKyM�T��IgF	�5)�����O}���2_BUF�F 2��� �p�2O�_�2��6_ M�R_d_�_�_�_�_�_ �_�_�_o3o*o<oNo�`o�o�o�o�o���ADCS ������ �L�O��+=Oa��dIO 2��kc +����� �������*� :�L�^�r��������� ʏ܏���$�6�J�~uuER_ITM��d������ǟٟ��� �!�3�E�W�i�{��� ����ïկ�����7Nx�SEVD��t�TYP����s���8���)RSTe�e�SCRN_FL +2��}���π�/�A�S�e�wϨ�T�P{��b��=NG�NAM��E��dU�PSf0GI��2�����_LOADދ�G %��%�DROP_�EI�TO_3�ϑ�MA?XUALRMb2��@���
K���_PR��2  �3�AK�Ci0��qO=_'X��Ӭ�P 2��;� �*V	����
* ���4��*�� '�`�	xN��z��� ���������1�C�&� g�R���n��������� ��	��?*cF X������� ;0q\� ������/� /I/4/m/X/�/�/�/ �/�/�/�/�/!??E? 0?i?{?^?�?�?�?�? �?�?�?OOAOSO6OpwObO�OD�DBG*� ��գѢѤO�@�_LDXDISA�����ssMEMO_{AP��E ?��
 �Ax$_6_�H_Z_l_~_�_�_K�F�RQ_CFG �����CA w@i��S�@<��d%�\�o�_�P�Ґ�����*Z`/\b **:eb�DXo jho�F�o�o�o�o�o �o;�O��dZ�`U�y|��z,(9 �Mt���1��B� g�N���r���������̏	���?�A�IS�C 1���K` � �O�����O���O֟�����K�]�_MSTR� �3��SCD 1�]��l�� ��{�����دïկ� ��2��V�A�z�e��� ����Կ������� @�+�=�v�aϚυϾ� ����������<�'� `�K߄�oߨߓߥ��� �����&��J�5�Z� ��k���������� ����F�1�j�U��� y��������������0T?x�MK��Q�,��Q�$M�LTARM�R�:?g� ~s�@����@METPU��@l��4�ND�SP_ADCOLx�@!CMNT7 *FNSW(FSTLIxi%� �,����Q�|�*POSCF�=bPRPMV��ST51�,� 4�R#�
g!|qg% w/�'c/�/�/�/�/�/ �/?�/?G?)?;?}? _?q?�?�?�?�?�1*�SING_CHK�  {$MODA�S�e���#E�DEV 	�J	�MC:WLHSI�ZE�Ml �#ETA�SK %�J%$�12345678�9 �O�E!GTRI�G 1�,� l �Eo#_�y_S_�}�F�YP�A�u9D"CE�M_INF 1��?k`)AT?&FV0E0X_�]�)�QE0V1&�A3&B1&D2�&S0&C1S0}=�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_�_o �3o��o���o� �"�4��X��� ASe֏���C� 0���f�!���q��� ��s�䟗�����͏>� �b���s���K���w� ��ٯ�ɟ۟L��� �#�����Y�ʿ�� ����$�߿H�/�l�~� 1���U�g�y����ϯ�  �2�i�V�	�z�5ߋ��ߗ���PONITO�R�G ?kK  � 	EXEC�1o�2�3�4��5��@�7�8
�9o��� ��(��4��@��L� ��X��d��p��|⪂�2��2��2��2���2��2��2��2���2��2��3��3��3(�#AR_GRP_SV 1��[� (�1@3>��?|�/�Q���6 `��@Q��>��zRM�A_D�sҔN��ION_D�B-@�1Ml  K�l yFH"b+��l FH��N �BL"FI-ud�1}E���)PL�_NAME !��E� �!De�fault Pe�rsonalit�y (from �FD)b*RR2��� 1�L�X�L�p�X  d�-?Qcu �������/ /)/;/M/_/q/�/�/�/f2)�/�/�/?�?,?>?P?b?t?f< �/�?�?�?�?�?�?
O�O.O@OROdOc	�6D�?�N
�O�OfP�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ �O�O2oDoVohozo�o �o�o�o�o�o�o
 .@o!ov��� ������*�<��N�`�r����� �Fs  GT��G�Me��x �ÏՍfd������ �(�6������
 �m�p~�h����� �� ����ğ֟�����:����
�]�m�f��	�`������į��:�oAb	����� A�  /� ��P����r������� ^�˿ݿȿ��%���R�� 1��	X ���, � ���� a� @D� M t�?�z�`�?f <|�fA/��t�{	ު�;�	l��	 ��x�J������ �� ��<�@���� ���·�K�K� ��K=*�J����J���J9��
�ԏC����t�@{S�\��(Ehє��.���I����>����T;f�ґ��$��3��´  �@��>�Թ�$��  >�����{�Uf��x`���� �
��������� �  _{  @T�����P �H �l�ϊ��-�	'� � ���I� � � �<�+�:������È=��ͨ��0Ӂ��N �[��n @���f���f�k���,�av�  '������@2��@�0�@�Ш���C��C>b C��\C����z��G�@��I����� )�Bb �$/�!��L��Dz �o�ߓ~��0���( �� -��������!���D�  |��恀?�ffG�*<� }�q�"1�8����>��bp$��(�(���P��	�������>�?����x���W�<
6�b<߈;܍��<�ê<���<�^��I/��A�{��fÌ�,��?fff?_�?&�� T�@�.�"��J<?�\��"N\�5���!��(�|� �/z��/j'��[0?? T???x?c?�?�?�?�?0�?�?5��%F��? 2O�?VO�/wO�)IO�O�EHG@ G@0~��G�� G}� �O�O�O_	_B_-_f_�Q_BL��B[�A w_[_�_b��_�[�_�� mO3o�OZo�_~o�o�o<�o���b��PV( @|po	lo-*cU�ߡA���r5�eCP�Lo�}?����#��5���W�s��6�Cv�q�CH3� j�t�����q�����|^(�hA� �ALf�fA]��?�$��?��;�°�u�æ�)�	�ff��C�#s�
���g\)�"��33C�
�����<�؎�G�B������L�B�s�����	";�H��ۚG��!G���WIYE���C�+�8��I۪I�5��HgMG�3�E��RC�j=�x�
�pI����G��fIV=�?E<YD�C<� ݟȟ����7�"�[� F��j�������ٯį ���!��E�0�i�T� f�����ÿ���ҿ� ���A�,�e�Pω�t� �Ϙ��ϼ������+� �O�:�s�^߃ߩߔ� �߸������ �9�$� 6�o�Z��~����� �������5� �Y�D� }�h����������������
C.(䁳3��/"���<���t��q3ǭ8����q4M�gu���q�Vw�Q�
4p�+4�]$$dR�Pv���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/�/X�/�/�/  %��/ �/+??O?:?s?/�_0�?�?�?�;�?�?@O�? OFO4O�rLO�^O�O�O�O�O�O�J � 2 Fs�wGwT�V�M�uaBO�|r�pp�C��S@�R_�to}_�_f_��_�|\!�W����_oo(o�z?̯��@@�z�DR�p�pk1�p�~
 6o�o�o�o�o �o�o);M_pq�ڊsa �����D��$MR�_CABLE 2}�� ]�J�T�LaMa?�PXMaLb�p�Z��&P��C�p�!O4>��B����!Y�4� �!E�h\��&��v�l  ���&P�v�wdN�{u0��$s8ca��F�� 6�H�eXT��6P� C$��Č��n��u	� 'z�"������� ��&P��C\���=��������� )z��~։��s9��T�,� >���b�������Ɵ�� Ο3�.��P�(�:��� ^���j��#� ���� ��;h�H�Z�l�;hw*��** �s�OM ��y����B�"���%�% 234567O8901ɿ۵ ƿH���� �� AQ� ��!
�z�n�ot sent 앺�W�T�ESTFECSA�LG� eg;jAQdȎ�ga%�
���@���$�r�̹�������� 9UD1:�\mainten�ances.xm�S�.�@�vj�DEFAULT�\~�rGRP 2���/  p� �J�%�  �%1st� mechani�cal chec�k��!���������E��Z�(��:�L�^��"��controller�����߰��D�����0 ��$�s�M��L��""8b���v��B�����������/�AC}�a�6����@dv���s�C���ge��. battery�&��E	S(:L^p�	�|�duiz�abl�et  D�а�R���/�"/4/s��gre�as��'f�r#-� |!�/�E��/�/��/�/�/s�
�oi0,�g/y/�/�/t? �?�?�?�?s��
�XֈW��1<X�AO�E
c?8OJO\OnO�OB�t��?O��'O��O_ _2_D_s�O?verhauE��L��R xXЌQ�_���O�_�_�_�_o�X�$�_0o����_o  �_�o�o�o�o�oo�o ?oQocoJ\n� ��o�)�� "�4�F���|��k� �ď֏����[�0� B���f����������� ҟ!���E�W�,�{�P� b�t�����矼��� �A��(�:�L�^��� ��ѯ㯸��ܿ� � �$�s�Hϗ���~�Ϳ �ϴ�������9��]� o�Dߓ�h�zߌߞ߰� ����#�5�G���.�@� R�d�v��ߚ������ ������*�y���`� ��O������������ ?�&u�J��n� ����); _4FXj|�� ��%�//0/ B/�f/���/��/ �/�/�/?W/,?{/�/ b?�/�?�?�?�?�?? �?A?S?(Ow?LO^OpO �O�O�?�OOO+O�O _$_6_H_Z_�O~_�O �O�O�_�_�_�_o o�P�R	 T"oOoao so�_�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z��������ԏ���
�� � ��Q?�  @�a �oW�i��{��fC�����̟aX;*�** �Q�V ��� �2�D��h�z��������_�S� �����կ7�I�[� ����ɯ/���ǿٿ#� ��!�3�}�����{� �ϟ��s�������C� U�g��S�e�w�9ߛߠ�߿�	�߉e�a��$MR_HIST� 2��U�� �
 \jR$ 23�45678901P*�2����)�9c_ ���R��a_����� ����=�O�a��*�x� ����r������� 9��]o&�J� ����#�G��k}4��d�S�KCFMAP  ]�U������`��ON�REL  �����лEXCFENB'
��!�FNC$/$JOG_OVLIM'd�\m �KEY'p%=y%_PAN(�"\�"�RUN`,p%��SFSPDT�YPD(%�SIG�N/$T1MOT�b/!�_CE_�GRP 1��U�"�:`��n?�c[? �?�؆?�?~?�?�?�? !O�?EO�?:O{O2O�O �OhO�O�O�O_�O/_ �O(_e__�_�_�_�_�v_�_�_�_o�׻Q?Z_EDIT4���#TCOM_CF/G 1��'%to�o�o 
Ua_AR�C_!"��O)T_MN_MODE6{�Lj_SPL�o�2&UAP_CPL��o3$NOCHEC�K ?� � Rdv�� �������*��<�N�`��NO_WAIT_L 7Jg50NT]a���UZ���_ERR?12	���ф��	��-�@���R�d����`O��}��| ��0
a�B����o����C��������,rV<� �� ?�U�ϟj����قPAR�AMႳ���N�oR�=��o��� = e������گ �ȯ��"�4��X�j�F�<�蜿��A�ҿ~�"ODRDSP�c�6/(OFFSET�_CAR@`�o�DsIS��S_A�`�ARK7KiOPE?N_FILE4�1��aKf�`OPTIO�N_IO�/�!��M_PRG %��%$*����h�WO�T��E7O�p���Z��  �'  Z"�÷"�G	 �V"�Z����RG_DS�BL  ���ˊ���RIENTkTO ZC����A(��U�`IM�_D���O��V~�LCT ����Gbԛa�Zd��_�PEX�`7�*�RA-T�g d/%*���UP ���{��������������/$PAL�������_POS_CHU��7����2>3�L��XL�p��$�ÿU�g�y��� ������������	 -?Qcu����Y2C���" 4FXj|�� ���� //$/6/@H/Z/l/~/�Y�� �.��/�/ςP�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO�/ �/LO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_)O;O�_�_�_�_�_ �_�_o o2oDoVoho�zo�o�o�_<���o�m ���~ BPw�m�m���~�jw8��w���� ��2�T��p��w���H��t	`���̏ޏ��:�o������ �2��pA�   I��j�`������ ���џ���@���#�)�Or�1�3���3� 8�>��, �\Ԡ�~� @D�  ��?���~�?� ���!�D������%G� � ;�	l��	 ��x�J젌����� ��<� ��� ���2�H(��H�3k7HSM5G��22G���GN�3%�R��oR�d��2�Cf��a��{���������/��3��-¸��4��>����𚿬���3�A�q�½{q�!ª��ֱ� "�(«�p=�2����� ��_{  @�Њ��_�  ��Њ��2���.�	'� �� ��I� ��  �V�,�=�������˖ß���  �y��n @"��]�<߼+"������-�N�Д߇  '�Ь�w�ӰC>��C��\C߰���Ϲ��ߤ!���@%�4���/��2�~�B��B�I�;�)�j客z+���쿱����������( �� -��#�������!�]�9�|�  q�?�ffaH�Z��� ������"��8� ����>�|P$��}�(� ��P��������\�?���� x� ���<
6�b<߈;܍��<�ê<���<�^�*�gv�A)ۙ�脣��F��?fff?}�?&�� ��@�.���J<?�\��N\��)������� ����ޤy�N9 r]������ �/&/�J/5/n/��	g/�/c(G@� G@0i�G�� G}���/??<?�'?`?K?�?o?BL
i�B��A�?y?�?|� �?K�?ů�/QO�/xO��?�O�O�O�Om��bs��n�t @|�O '_�OK_6_H_�_lS��!A��RS�i�Cn_�_xj_0O�]?��o�oAo,o¹�Wi����ToC���`CH�Qo>Jd�`a�a@�Iܚ>(hA�� �ALffA�]��?�$�?����ź°u��æ�)�	ff���C�#�
ܢopg\)��3�3C�
������<��nG��B���L��B�s�����	0źH����G��!G���WIYE����C�+�½I�۪I�5�H�gMG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo�� �
��U�@�y�d��� ������я����� ?�*�c�N���r����� ���̟��)��9� _�J���n�����˯�� �گ�%��I�4�m� X���|���ǿ���ֿ ���3��W�B�Tύ� xϱϜ���������	� /��S�>�w�bߛ߆� �ߪ߼�������=��(�a�L�(q���)����Z�������a3�8�������a4Mgux�����a�VwQ��(�4p�+4�]B�B���p�����������UPbP���Q O%x�1[FjR�������  C���I 4mX�8
O������.//>/d/R/�Rj/|/�/�/�/�/�/:  2� Fs�gGT]�&6�M�eBmpX�R�P�aC��3@�_ p?�?�?�?�?�?�=�S�OO)O;OMO�c�?���@@�jJ��`�`�1�`�^
 TO�O�O �O�O�O_#_5_G_Y_�k_}_�_�_�j�A �����D��$�PARAM_ME�NU ?B���  �DEFPULS�E{	WAIT�TMOUTkR�CVo SH�ELL_WRK.�$CUR_STY�L`DlOPT�Z1ZoPTBooibC�?oR_DECSN `���l�o�o�o &OJ\n������QSSREL_ID  >��
1��uUSE_P�ROG %�Z%8�@��sCCR` ��
1�SS�_HOST7 !�Z!X����M�T _���x�������L�_TIME�b �h��PGDE�BUG�p�[�sGI�NP_FLMSK��E�T� V�G�PG�Ar� 5��?��CyHS�D�TYPE�\�0��
�3�.� @�R�{�v�����ï�� Я����*�S�N� `�r����������޿ ��+�&�8�J�s�n���ϒϻ�G�WORD� ?	�[
 	�PR2��MA9I�`�SU�a��cTEԀ���	Sd�COL��C߸��L� C�~��h�d*�TRACE�CTL 1�B���Q ��m n'��0�ށ�_DT Q�B������D � ���q����
�����1�@� �@⨐�@�@�U � �	����U�������&�U�.�������U���&��.��6�U�>��F�
H�H�H����������K H� ������5��������U�������&��.��6��>�U�g��y���G�������Ѯ��� ���� ��������/�A�S� e�w��������������������O
��OO�Ug��X��XXX
X�Xf�����V�V�V�V���V��V��V��V���V��V��V���!�������@�� �� 2DNhz �f����-�?� ���?�?�?�������� ��d5(O:OLO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�P�$Or������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~�f���� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo��o�o�o�o�o�a�$�PGTRACEL�EN  �a  ���`���f_UP �/���q'pq� p�a_CFG7 �u	s�a p�LtLtfqw|pqz  �qu�4rDEFSPD ��?|�ap���`H_CONFI�G �us U�`�`d�t��b �a�qP�t�q���`��`IN7pT�RL �?}_q8l�u�PE�u��w�qLt�qqv�`WLID8s�?}	v��LLB 1��y� ��B�pB94Ńqv �އ�؏	�s << �a?��'�� �A�o�U�w������� ۟��ӟ��#�	�+�Y�v�񂍯����ï
���������/�u�GRoP 1ƪ��a�@�j��hs��aA�
D��� D@� Cŀ7 @�٭^�t�q0�����q�p���.� ���Ⱦ´���ʻB�)�	���?�)��c��a>��>��,��Ϻ��ζ� =49X=H�9�� 
����@�+�d�O����s߬�o߼�����  #Dz���`
��8� ��H�n�Y��}��� ����������4��X��C�|���)��
V�7.10beta�1Xv A������!�����?�!G�>\=�y�#��{33A!��@��͵���8wA��@_� A�s�@Ls���� ��"4FX�LsApLry�ā�_��@l�ͯ@�33q�`s���k��Anff��a��ھ��o)�x�� �a r�T�n�t�����	t�KNOW_M�  |uGvz�SV7 ��z�r� &����>/�/PG/�a��y�MM���{� ���	^u (l+/�/',_t�@XLs	����@���%�"�4�.N�z�MRM��|-TU�y�c?u;e�OADBANFW�D~x�STM�1 �1�y�4Garra_B�2Sem��?~s�;Co�2��O�7��3Antena�_Full @� �VODe�qH��^OpO �O�O�O�O�O�O!_ _ _W_6_H_�_l_~_�_��b�72�<�!4�_ � �<�_�_N�3 �_�_
oo�749oKo]ooo�75�o�o�o�o��76�o�o�77 2DVh�78��X���7MA�0���swwOVLD � �{�/a�2P�ARNUM  p�;]��u�SCH*� 8�
����ω�3�UPD��[�ܵ+�>wu_CMP_r -���0�'�5C�ER�_CHKQ���`�1�"e�N�`�RS>0��?G�_MO�?_���#u_RES_G
�0��{
Ϳ@�3� d�W���{�������� կ���*�����P��O��8`l��� ����`��ʿϿ��` �	���1p)�H�M� ��phχό���p��x�����V 1��5|�1�!@`y�ŒTHR_INR>0�/�Z"�5d:�MASmSG� Z[�MNF��y�MON_QUEUE ��5�6ӐV~  #tNH�U��qN�ֲ���END�����EXE������BE������OPT�IO������PROGRAM %���%��߰���TA�SK_I,�>�OCFG ά�]���^��DATAu#�����Ӑ2�%B�T� f�x���5��������������,>P�IWNFOu#� ���� ����� '9K]o��� �����/lx�� � ;���ȀK�_�����S&ECNB-�b-&q�&2�/ڝ(G��2�b+ �X,		��=�{���/��@��P4$�0��99)�N'�_EDIT ����W?i?��WERF�L�-ӱ3RGAD�J �F:A�  �5?Ӑ�5Wј6���]!֐��??�  Bz�WӐ<1Ӑ�%�%O�8�;��50!2��7�	�H��l0�,�B=P�0�@�0�M�*�@/�B *�*:�B�O�F�O2��D��A�ЎO�@O	_�,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_�_o �_o�_�_
o�o.o�o jodovo�o�o�o�o�o �o\XB<N� r����4��0� ��&���J������� ����������x� "�t�^�X�j�䟎��� ʟğ֟P���L�6�0� B���f���������(� ү$������>��� z�t��� Ϫ����� �l��h�R�L�^�DX�	���ώ0�� ���t$ :�L��o�
���ߥ��7PREF S��:�0�0
�5?IORITYX�M6}��1MPDSPV��:
B �UT��C�6�ODUCT���F:��NFOG[@_�TG�0��J:?�HI?BIT_DO�8���TOENT 1��F; (!AF�_INE*������!tcp����!ud��8�!�icm'��N?�X�Y�3�F<��1)�� �A�����0� ����������'  ]D�h�������*>��3���9
BOTf�3>�)��2�B�G/�LC���4�;LFJAB,  ���F!/�/%/7/�5�F�Z@�w/�/�/�/�3&�ENHANCE S�2FBAH+d�?�%;�������Ӓ1��1PORT_N�UM+��0����1_CARTRE�@��q�SKSTyA*��SLGS�������C�U�nothing�?�?OO�۶0TEMP �N�"O�E��0_a_seiban|߅OxߕO�O �O�O�O_�O'__K_ 6_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1U@e� v����������Q�<�u�.IVE�RSI	�L��� �disabl�e�.GSAVE ��N�	267_0H771|�h���!�/��9�:� !	^�4�ϐ����e��͟ߟ������9�D�C-Å_y� +1���������ő����Ǻ�URG�E� B��r�WF Ϡ��-��9�W�����l:WRUP_DELAY �=�n�WR_HOT �%��7��/p��R_NORMALO��V�_�����SEMI𓿹�����QSKI%Po��97��xf�=� b�a�sυ�H��ʹ��� ���������&��J� \�n�4�Fߤߒ����� �߲���� �F�X�j� 0��|�������� ���0�B�T��x�f����������ãRBT�IF�5���CVT�MOU�7�5����DCRo���� �T�A�:�CC�avC��>�;P>�[�a:�_�H�� ��c��^���?�S�`kϻ�4�HϘ�� �<
6b<߈�;܍�>u.��>*��<��� �P0���2 DVhz��������,GRDIO�_TYPE  �v��/ED� T_?CFG ��-BH]�EP)�2���+ ��B� u �/�*��/�?�/ %?=�/V?�}?�Ϟ? ���?�?�?�?�?O
O @O*Gl?qO��8O�O�O �O�O�O�O�O�O_<_ ^Oc_�O�__�_�_�_ �_�_o�_&oH_Mol_ o�oo�o�o�o�o�o �o�o"DoIho* j������� .3�E��f� ���x� �������ҏ�*�/� N��b�P���t����� Ο��ޟ�:�+���R'?INT 2�R��!=�1G;� i�{���"���8f�0  ��ӫ������ M�;�q�W�������˿ ���տ�%��I�7� m��eϣϑ��ϵ��� ����!��E�3�i�{� aߟߍ��߱����������A���EFPO�S1 1�!)  x���n#�� �����������/� �S���w����6��� ��l�������=O ����6���V� z� 9�]� ���Rd�� �#/�G/�k//h/ �/</�/`/�/�/?? �/�/?g?R?�?&?�? J?�?n?�?	O�?-O�? QO�?uO�O"O4OnO�O �O�O�O_�O;_�O8_ q__�_0_�_T_�_�_ �_�_�_7o"o[o�_o o�o>o�o�oto�o�o !�oEW�o>� ��^����� A��e� ���$����� Z�l�����+�ƏO� �s��p���D�͟h� 񟌟�'�ԟ�o� Z���.���R�ۯv�د ���5�ЯY���}��� *�<�v�׿¿����π��C�޿@�y��e�2 1�q��-�g��� ��	��-���Q���N� ��"߫�F���j��ߎ� �߲���M�8�q��� 0��T�������� 7���[�����T��� ����t�����!�� W��{�:�^ p��A�e  �$��Z�~ /�+/���$/�/ p/�/D/�/h/�/�/�/ '?�/K?�/o?
?�?.? @?R?�?�?�?O�?5O �?YO�?VO�O*O�ONO �OrO�O�O�O�O�OU_ @_y__�_8_�_\_�_ �_�_o�_?o�_co�_ o"o\o�o�o�o|o �o)�o&_�o� �B�fx��%� �I��m����,��� Ǐb�돆����3�Ώ ���,���x���L�՟ p�������/�ʟS���w�����ϓ�3 1��H�Z������6� <�Z���~��{���O� ؿs����� ϻ�Ϳ߿ �z�eϞ�9���]��� ����߷�@���d��� ��#�5�G߁������ ��*���N���K��� ��C���g������ ��J�5�n�	���-��� Q���������4�� X��Q��� q���T� x�7�[m �//>/�b/��/ !/�/�/W/�/{/?�/ (?�/�/�/!?�?m?�? A?�?e?�?�?�?$O�? HO�?lOO�O+O=OOO �O�O�O_�O2_�OV_ �OS_�_'_�_K_�_o_ �_�_�_�_�_Ro=ovo o�o5o�oYo�o�o�o �o<�o`�o Y���y��&� �#�\�������?�xȏ����4 1�˯ u�����?�*�c�i��� "���F����|���� )�ğM�����F��� ��˯f�﯊����� I��m����,���P� b�t������3�οW� �{��xϱ�L���p� �ϔ�߸������w� bߛ�6߿�Z���~��� ��=���a��߅� � 2�D�~��������'� ��K���H������@� ��d�����������G 2k�*�N� ���1�U� N���n� �/�/Q/�u// �/4/�/X/j/|/�/? ?;?�/_?�/�??�? �?T?�?x?O�?%O�? �?�?OOjO�O>O�O bO�O�O�O!_�OE_�O i__�_(_:_L_�_�_ �_o�_/o�_So�_Po �o$o�oHo�olo�oۏ�5 1����o�o �olW��o�O� s���2��V�� z��'�9�s�ԏ���� �����@�ۏ=�v�� ��5���Y��}����� ۟<�'�`�������� C���ޯy����&��� J����	�C�����ȿ c�쿇�ϫ��F�� j�ώ�)ϲ�M�_�q� �����0���T���x� �u߮�I���m��ߑ� �������t�_�� 3��W���{������ :���^�����/�A� {����� ��$��H ��E~�=�a �����D/h �'�K��� 
/�./�R/��/ K/�/�/�/k/�/�/? �/?N?�/r??�?1? �?U?g?y?�?O�?8O �?\O�?�OO}O�OQO��OuO�O�O"_t6 1�%�O�O_�_ �_�_�O�_|_o�_o ;o�__o�_�oo�oBo Tofo�o�o%�oI �omj�>�b �������i� T���(���L�Տp�ҏ ���/�ʏS��w�� $�6�p�џ������� ��=�؟:�s����2� ��V�߯z�����د9� $�]��������@��� ۿv�����#Ͼ�G�� ���@ϡό���`��� ��ߨ�
�C���g�� ��&߯�J�\�nߨ�	� ��-���Q���u��r� ��F���j������� �����q�\���0��� T���x�����7�� [��,>x� ���!�E�B {�:�^�� ���A/,/e/ /�/ $/�/H/�/�/~/?�/�+?�/O?5_GT7 1�R_�/?H?�?�?�? �/O�?2O�?/OhOO �O'O�OKO�OoO�O�O �O.__R_�Ov__�_ 5_�_�_k_�_�_o�_ <o�_�_�_5o�o�o�o Uo�oyo�o�o8�o \�o��?Qc ���"��F��j� �g���;�ď_�菃� �����ˏ�f�Q��� %���I�ҟm�ϟ��� ,�ǟP��t��!�3� m�ί��򯍯���:� կ7�p����/���S� ܿw�����տ6�!�Z� ��~�Ϣ�=ϟ���s� �ϗ� ߻�D������ =ߞ߉���]��߁�
� ���@���d��߈�#� ��G�Y�k�����*� ��N���r��o���C� ��g����������� nY�-�Q� u��4�X�x|b?t48 1�? );u��/;/ �_/�\/�/0/�/T/ �/x/?�/�/�/�/[? F???�?>?�?b?�? �?�?!O�?EO�?iOO O(ObO�O�O�O�O_ �O/_�O,_e_ _�_$_ �_H_�_l_~_�_�_+o oOo�_soo�o2o�o �oho�o�o�o9�o �o�o2�~�R� v���5��Y�� }����<�N�`����� ����C�ޏg��d� ��8���\�埀�	��� ��ȟ�c�N���"��� F�ϯj�̯���)�į M��q���0�j�˿ ��ￊ�Ϯ�7�ҿ4� m�ϑ�,ϵ�P���t� �Ϙ���3��W���{� ߟ�:ߜ���p��ߔ� ��A����� �:�� ���Z���~����� =���a���� ������MASK 1���������XNO  ���� ?MOTE  ��R_CFG ��Y����PL_RGANGUP���OWER ���� �A��*S�YSTEM*P�V9.3044 ��1/9/2020� A � ����RESTART�_T   , �$FLAG� �$DSB_SIG�NAL� $U�P_CND4P���RS232r� � $COM�MENT �$DEVICEU�SE4PEEC$�PARITY4O�PBITS4FL�OWCONTRO~3TIMEOUe�6CU�M4AU�XT��5INTE�RFACsTATeU�JCH� t $O�LD_yC_SW� 'FREEF?ROMSIZ ��ARGET_DI�R 	$UP?DT_MAP"� TSK_ENB"�EXP:*#!jF�AUL EV!�RV_DATA��  $n E��   	$VA�LU�! 	j&G�RP_  � {!A  2� �SCR�	� �$ITP�_�" $NU�M� OUP� �#T�OT_AX��#D�SP�&JOGLI��FINE_PC�d�OND�%$�UM�K5 _M�IR1!4PP TN�?8APL"G0_EXb0<$�!� 814�!{PGw6BRKH��;&NC� IS :�  �2TYP� �2��"P+ Ds�#;0B�SOC�&R N�5DUMMY164�"�SV_CODE_�OP�SFSPD__OVRD�2^�LDB3ORGT-P; LEFF�0<G�� OV5SFTJR3UNWC!SFpF5�%3UFRA�JTO~�LCHDLY7RECOVD'� �WS* �0�E0RO��10_p@  � @��S NVwERT"OFS�@9C� "FWD8A�D<4A�1ENABZ6�0�TR3$1_`1F�DO[6MB_CM��!FPB� BL_MP��!2hRnQ2xCV� "' } �#PBGiW|8AMz3\P��U�B�__M�P�M� �1�AOT$CA� �PD�2�PHBK+!:&a�IO�4 eIDX+bPPAj?a$i�Od7e�U7a�CDVC_DBG"�a;!&�`�B5�e1�j�S�ey3�f�@ATIO� ���AU�c� �S&�AB
0Y.#0 �D��X!� _�:&?SUBCPU%0SIN_RS�T, �1N|�S�T!�1$HW_C1�"]q.`<�v�Q$AT! � ��$UNIT�4|�p�pATTRI= ��r0CYCL3N�ECA�bL3FLT?R_2_FI9a7��c,!LP;CH�K_�SCT>3F�_�wF_�|8��zFqS+�R�rCHAGp��y��R�x�RSD��@'�1E#&7`_T��XPRO�`@S�E�MPER_0�3T�f�]p� f��P�D�IAG;%RAIL�AC�c4rM� LOh�0�A�65�"PS�"b�2 -`�e�SPR�`MS.  �W�Ctazf	�CFUNC�2��RINS_T�.!(�w��� S_� �0�P�� 	d���WARL0bCBL'CUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!2��8�3�TID�S���!� $CE_R�IA !5AFDpPbC~��@��T2 �1C9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@H�RDYOL1	PRG�8�H��>1(�ҥM�ULSE =#Sw3.��$JJJ6BKG�FKFAN_ALMsLV3R�WRNY��HARD�0+&_P� "��2Q���!�5_,�@:&AU�Rk��?TO_SBRvb���� ƺ�pvc�޳MPINF�@�q�)�N��REG'd~0V) x0R�C�1DAL_ �\2FL�u�2$M@Ԑ(�#S��P� `�6g�CMt`NF�qsONIP�qEIPP� 9a$Y���!�"�!o� �o3EGP��#@��AR� �c�5�2�����|5AXE��'ROB�*RED&�&WR�@�1_=��3CSY�0ѥ0_�Si��WRI�@�ƅpST��#��0*@� �q	���3��� B� �A�ֺ3�D�POTO�� �@ARY�#��!���d�!1FI�0��$LINK��GT5H�B T_���A���6�"/�XYZt+"9�7G�OFF�@R�.�"���B� �l����A3$ ��F�I�p���4�4l��$_Jd�"(B�,a������8�"q����d��Ck6DUR���94�TURT�XZ�N����Xx��P��FL/�@s��l�P���30�"Q 1�� K
0M:$�53�]q7�SuD�Sw#ORQɆ�!�����Q7��0O[�ND�=#�!#�N1OVE8��M� ��R��R��Q!`P.!P! OAN}q 	�R����990� �b rJ9V����v��!ER1��	8�E��@n D�A��p��嘕Ă���v�AX�C�"��`�q�s ���0~3�~ F�~e�~�~E�~1��~Ҡ{Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�Ҡ��Ҡ�Ҡ�!)D7EBU}s$x���0삼!R*�AB�a�8A2V`|r 
 �"�c���%�Q7�7 �173�7F�7e�7 �7E�������LAB����yp�cGGRO�p��}��PB_ҁ ��̓��ð��6�1���5���6AND��8p�a3���-G �Q����AH�PH��p2�NTd��Cs@V�EL؁�}A��F��SERVEs@��� $����A!�!�@POR}�KP�иA� �B���	��]$�BTRQ�
�CdH��@
�G��2	�E�b��_  l8b��Q�ERR��R�I�P�@�FQTOQ�� L�}��YVĀeG�E%�\��C�RE�  ,h�A�EP
�RA�Q? 2 d�R7c��D�A ���$F ׂ��m���BO�C��P  �8[COUNT�� �,�SFZN�_CFG�A 4�p%��rT\zs�a�#�`pJp�R�Q(a�� �� MGp+����`0�OGp�eFAq����cX8еk�ioQ��$'ѴDp8�Pz����HELA�-b� 5��B_BA�S\RSR$�`�"2�S��L�!p1�W!pU2Dz3Dz4Dz5Dz�6Dz7Dz8�WqR�OO���P�1�NL��� �AB�C
�"pA[CK�&IN�PT+��W�U��	�k��y_P�U8�~�|�OU�CP���%�s�Vl���YT�PFWD_KAR�KQ-�:PRE�D�P8����QUE$�Ā 9 )���~���IU��#�s/���@�/�SE�M1ǆ1�A�aS�TY�tSO����D�I�q��Qc��X��_�TM9�MANRQ� �/�END��$�KEYSWITCaH2�G����HE)��BEATMz�PE���LEJR���0x�U�F�F��G�S�DO/_HOM��Oz��pEFPR��SbJ����uC��O��7P�Q�OV_M��}�c�IGOCM���1�BvsHK�� D,�$&�a`U2R��M��a��r +�FORC*�WcAR�.� uOM��  @�$�㰰U��P�1��g���U3��4��S�POW��Lz��R%�UNLiO�0T�ED��  �SNP���S.b 0N�AD�Da`z�$SIZ�*�$VA�0�UM_ULTIP�r����Az� � �$��ƒ���S�Qc�1CFPv�FRI	Fr�PSw���ʔf�{NF#�ODBUxЀR@w������F��:�I�Ah����������S|"p�� �  ��cRTE���SG%L.�T�x�&C`G�x�3a�/�STMT��2`�P����BW9 0��SHOWh�qBANt�TPo���E�Ц����@V_Gvsb �$PC�0X�PoFBv�P�ȋSP��A�p���`V�D��rb� �+QA002D.ҝ��6ק�6ױ�6׻�6�5�4�64�74�84�9
4�A4�B4و�6ׇ17�}�6�F4� ��@�@����Z����t�1��U1��1��1��1��U1��1��1��1��U1��23�2@�2M�U2Z�2g�2t�2��U2��2��2��2��U2��2��2��2�م2��33����M�3�Z�3g�3t�3��3���3��3��3��3���3��3��3��3���43�4@�4M�4�Z�4g�4t�4��4���4��4��4��4���4��4��4��4���53�5@�5M�5�Z�5g�5t�5��5���5��5��5��5���5��5��5��5���63�6@�6M�6�Z�6g�6t�6��6���6��6��6��6���6��6��6��6���73�7@�7M�7�Z�7g�7t�7��7���7��7��7��7���7��7��7��7����VPv�U�BG �@�09r
��|���A x �0YR���  �BM�@�RP�`�4Q_�PR��@[U�AR��DSMC4��E2F_U��=A���YSL�P�@ �  �ֲ>g���ଐ��iD��VALAU>e�pL�A�HFZA�ID_L���EHI��JIh�$FILE1_ ��D�d$Ǔ��XCSA�Q h��0!PE_BLCK�z�.RI�7XD_CPUGY!�GY�Ic�O
T��PY.��R ? � PW`�pl���QLAn�S�Q��S�Q�TRUN_FLG�U�T�Q�TJ��U�Q�T�Q�UH��T`~�T	 �T2L��_LIz�  ]�pG_OT��P_EDIU��T2�`7c ?bة�p�BQh�)a�TBC2 �! �%�>��P��a�7aFTτ�d݃TDC�PA�N`�`aM�0�f�a�gTH��"U��d�3�gR�q�9�ERVEЃt݃�t	��a�p�` �"X -$EqL�ENЃRt݃Ep�pR1Av��Y@W_AtSi1Eq�D2�wMO?Q�S���pI�.B�A0�y�4Ep�{DE�u���LACE �CCC8�.B��_MA��v8��w�TCV�:��wT,�;�Z�P���sP�~��s�J�AՉM����J���uā�uQq2ѐ����݁�s�JK��VK@������	���J��l��JJ�JJ�AAL�<��<�6�d�:�5�cm�N1a�Pm�,��DL�p_\�nŰ���aCF
��# `�0GROUP�@J�Բ��N�`C^�~ȐREQUIRr�ÀEBUu�Aq��$T�p2"��Bp�8�a	��d$ \?@qhoAPPR��CLB�
$H`N;�CLOD}`K�S�e`��u
�a.I�% �3�M�`�8l��_MG񱥠�C �"P����&���B{RK��NOLD����RTMO6a�ޭ��J6`�P>��p���p��pZ��pc��p6�+�7+�<�   |@r�d&� ��lr��������PATH��������qx��䋠�%0A��SCA�ub��<���INDrU�C�p�q�C�UM�Y�psP����A� q/ʤ�/�E�/�PA�YLOA�J2L��0R_AN�ap�L��Pz�v�jɆ���R_?F2LSHRt��LO{�R�������ACRL_�q������b�d�H�@B$yH��"�FLEX>��.`BJ�f' P�(��o�o+�py�J>Du( :Qcv �p����fe��po��|F1���-�� ����]�E�� *�<�N�`�r�����4� Q�������A�c���ɏHۏ���T��2�X:A ��������� �)�;�?�H�6�Z�c��u������0?Ь�) ���`��˟ݟ�`�0A1TF�𑢀EL���a���J�(��JE�۠CTR��A�TN��1�HAND_�VBB>ѯ@�*� $��F2���dƝCSW��x���+� $$M�����0 ˡ�ڡ�������A�@g����A)��A(���@˪A٫A� ���`P˪D٫D�P2ȰG�P�)STͧ�!4ک�!N�DY�P9� ���#%��Fp���Ѫǀ��i����������P 3�<�E�N�W�`�i�r����, ��ԓ�� n�5m��1AS�YMص.@�ض+A������_`��	� ��D�&�8�J�\�n�Ju�&��ʧC�I��.S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R�� &T��3TWV�͢���&��ߪU��/�7�;�f�`HR`ta-���QQ�1�DI��Op�T���P��. ; 
*"IAA*���$aG��2C2cJ�$y�I��P �/ � �M�E�� Mb�R4AT�PPT�@� ��ua�����P�l@zh�a�iT��@�� $DU�MMY1E�$P�S_D�RF�u$�f3�FLA���YP���b}c$GLB_T��Uuu`�1����EQa0 �X(���ST�����SBR�PM21�_V��T$SV_�ER��O_@KscsC)LpKrA��O'b�P�GL�@EW��1 �4��a$Y|ZB|W�s怯��AN`���`�sU�u2 ��N�p�@$GI�U}$�q �1u�q�p��3 L����v^B}$F^BE^�vNEAR��NK�yF8���TANCK�ΩJOG��� �4H`$JOIN�T����x��qMSE]T��5  �wE��H�� S�����6��  MU��?����LOCK_F�O����PBGLV�HGL�TEST�_XM>���EMP�t����r̀$1U�Гr��22���sB,�3���Ҁ,�1Mq�CE���sM� $K�AR��M�STPD�RA�pj�a�VECX��{�e�IU,�41�{HEԀTOOL�ڠ�V�RE��IS�3����6N�A�AC)H���5��O�}cj�d3���pSI.��  @$RAI�L_BOXE���ppROBO��?�~pqHOWWAR*�x��`�ROLM�b B���S��
�5����O_F� !ppHOTML5�Q��h����RGU�CH���7m�I`R��O��8`m��v�z���OU��'9 tpp(�14AX�̀��PO֡%PIP��N��
��ڑS�,�����COR�DEDҀް̠5�X�T��q)"rP� O�4` : D pOBP!"Ҁ{�j��cpj�^@$SYS�j�ADR#�Pu`T�CH� ; ,���EN�RZ�Aف_��t״����PV�WVAPa< �� p��r�UPRE�V_RT]1$E�DIT�VSHW�R�7v;���q��@D_`#R�+$HEADoA�Pl��A$�KE�q�`C�PSPD��JMPz��L�U�TR��Fd=r�O�϶I�5S#CiNE��$�_TICK�AM�X��q��HN-q�> @t������_�GP��[�STYѲ�LOq�s��Ҫ��?�
�Gݵ%�$���t=7pS !$Q��da�e!`�f9P�0�SQUd� �<�b�ATERCy`|zuS�@ �p�Cp����d�%Oz`mcO�IZ�d�q�e�aPRM��a8�����PUQH�_DO�=�ְXS��K�VA�XIg�f�1�UR � ��$#�Е��� Y_����ET��Pۂ����5f�F�7g�A��!�1�d9�2�;�SR|Al�о���#�� 5��#��#�)#�) i�>'i�N'i�^&{��� �){����2��C�����C��WOiO{O�D�S}Cp B hppcDS(�k��`SP`&�ATL �I����¼bADDRESz��B'�SHIF��^"�_2CH#���I&p��TU&pI�� Cm�CUSSTO��ޡV��IbADȲ�c�0
��
ݢV�X�R`E 	\�����f�7��tC�#	���F��ir�t�TXSCRE�El�F�P��TICNA�s�p��t��8���0G T��fp �b��eqBp&uᦲu�$#�RRO'0R����}�!����UE��H# ��0���`S�q��'RSM�k�UV����V~!�PS_�s�&C �!�)�'C��Cǂz"�� 2G�UE©4Ibvr�&8�GMTjPLDQ��Rp�~z��BBL_�9W�`R`J �f�>25O�qJ2LE�U3x"�T4RIGH^3�BRDxt�CKG�R�`�5TW��7�1WIDTH�H�����|�a��P�UIu�sEY��QaK d�pЅ�A�J�
�4�BACCKH��b�5|qX`sFOD�GLABS��?(X`I�˂$�UR(�9@���0^`H>4! L 8�QR�!_k��\B_`R�p͂������HBO�R`M���w0Uj0�CRۂM�LUM�C��� GERV��p�0P<�j�4NV`��GE=B0#���]�t�LP�E��	E��Z)Wj'Xz�'XԐ&Y5$[6$[7$[8	R���3�<��ԾfԑŁS��M��1USR�tO �<��^`U�r�rF�O
�rPRI��mx����PTRIP�m�UNDO��P�p��`m�4��l��#���� qQWB�P7�G s�aTf�H�RbOS�a�gfR��:">c��.qR���s�~�b*��A$�UQ.qS�o�o�#R)�N>cOFF���pT� ��cOp 1Rh�t/tS�GU���P.q��JsETw�1S�UB*� f�E_�EXE��V��>cW]O>� U�`^gF��WA'��P�q!@=� V_DB�s�pN�BSRT�`
�VҘQ�r��OR��uRAU��tT�ͷ�q9_���W |%�͸�OWNA`޴$S#RCE � ��D��\��MPFIA�p��ESPD������C����Gƒ� +�5��!X# `�`�r޴��7COP�a$��C`�_w������rCT�3�q���qƒ�`���@� Y"SH�ADOW�ઓ@�_UNSCA��@��4�M�DGDߑ��EGSAC�,me�G�oZ (0NO�@��D<�PE�B��V�W� �G���![ 7� ��VEE#��ڒANG�$��c�|�cڒLIM_X�c ��c� ����#��0`� 퐾�VF� �sO�VCCjв�\ՒC{�RAlצ���.RpNFA��%�-E��Z`G� ^03[�C`DEĒ��� STEQ1���@� ꁻ@I��`+0����`8����P_A6�r����K��!]� 1Ҡ�����\����CPC�@]�DRIܐ\�͑V#Ѐ����D�TMY_UBY �T���c��F!���Y�1븲���P_V�y���LN�BMQ1$n��DEY��EX��e��MU��X�MƓ US�!���P_R�����P� ߖG��PACIr�ʐf�ᔟ�@�c�´c���#�EqB���a.2B����^S ܀GΐP�H���@C�R~``�_�0��@3!�1zr	�e�R�SW��p�00��S�6�O�Q�1A� X�#�ME�UE��00�`VC�HKJ�`�@p����U� �EAN��ٖp�pXն�C�MR�CV�!a ��@O*��M�pC�	��s����REF*7
��� �����/��P��@��� @��b��֗�_Y��� ���ۣ��Q$3���p���C��$b �����%���Q��$GROU� �c�����2ʠ]��I2^0��U` 0_�I,�o � ULա`��C�&�rAaB�?�NT ���������A���Q��K�L����õ��A���Q��T a$c tf�`MD�p8�HU����SA�CMPBE F  _�ARr�p@����XS	�qVGF/�b#d, &�@M�P^0۰UF_C !���z �ROh0"+���@���0C�UREB���3RI��
IN�p� ����d��d��ca��INE�H�y��0V@�a-�걗��W�������C��i�LO�}�z�@0�!�QNSI��݁���c$&x�c$&.�X_PE-�YW+Z_M�ڒWD�I�$�" �+R�'�rRSLre �$/�M
`�RE�C7�Gd�۰�̵ҭ� q����u��Ȑ�������S_P�VnP �_�VIA�vf� �~pHDR�p�pJO�P��_$Z_UP��a_LOW�5�1J�dA���LINubEP�?�tc_i�1�1���@��G1@�V�xg{ 5X�PATHP= X�CACH$��]E��yI�A��{�C�)�ID3FA�ETD��H��$HO�pO�b@�{�d6�F����<��p�PAGE�䁀�VP�°�(R_SI	Z��2TZ3�-X�0U̲q�MPRZ��IM5G���AD�Y��MRE��R7WGP���8�p��ASYN�BUF�VRTD��U�T7Q�LE_2�D-��U��`CҡU�1��Qu��UECCU��VEM��]EDb�GVIRC�Q�U�S��B�Q�LA��p�N�FOUN_�DIAuG�YRE�XYZ�cE�WѴh8�dpq2a`T��2�IM�a�V�|be��EGRABBr��Y�a�LERj��C4���FC-A�65�04x��7u��@G��h�'�`�CKLAS�_@l�BA��N@i  $G��T��� @ݲմq$BAƠwj �!q�eb��uTYSp�H����2��I�t:b�f���B)�EVE����PaK���fx��GI�p�NO��2�AB_H�O����k � @���
8�Pi�S�0�ޗ��RO�ACC�EL?0=���VR_�U7@�`��2�p��AR��PA��̎K�}D��REM_But3 ��#�JMX ��l�t�$SSC��U �"#���QN@m� � �S�P�N�S��LEX�vn =T�ENAB 2¼W@��FLDRߨF�I�P�t�ߨ(Ğ�ޱ��VP2HFo'� ��V
Q MV_PI��8T @󐉰�F@�Z�+�#��8�8�#��GAB���LO9O��JCBx��w�"SCON(P�PLCANۀ�Dp�3F�d�v�9PէM��Q ;����SM0E�ɥ�8�ɥWb72$`<�8T̸�,`RKh"ǁVAsNC���1R_Ou N@p (�-#<#cp��c2��R_A/�N@q 4������`p	�^����r hn�p��1^�&OFF`�|�p�`��`�DEA��
�P,`SK�DM�P6VIE��2q �w��@���rs <C {���4���r�{7��D�����C�UST�U��t� $G�TIT1�$PR\��OPyTap ��VSF��
�su�p�0`r&�,*���MOwvI�|��ĄJ�����eQ_$WB��wI���� @�O3�@�XVRx�xmr��T�� ��ZABC��y �op����)�
�Z�D$�CSCH��z Lu����`�2�%P0C ��7PGN ��x<��A��_FUNH���@r�ZIPw{,I��LV,SL��~��np�ZMPCF���|��E����X�DMY_LNH�=����M|��} �$�A� ]�CMCM�� C,SC&!��P~�� $J����DQ�������������_�Q,2����U�X�a\�UXEUL ��a������(�:�x(�J���FTFL���w��Z�~�?@+�6� ̐��Y�@Dp  8/ $R�PU��> �EIGH����?(��iֱ��0��et�� �a�����$B��0�0@�	�_SH�IFD3-�RVV`FL�@��	$5��C�0���&!������b
h�sx�uD�TRR��V̱��P� H���!� ,�������s �4A�RYP���%����?�%����"�%!� �H�(UN0���"�2 ����ёЌq0�GSPDak����P��O�����0��mp���"!NGVER`q �iw+I�_AIRPURG�E  i  �i/�F`E�Tb� ��+  � h2I�SOLC  �,"�"�!���!�%�²P+�_/*OB��D�m�?@�!�H771   34n?�?�9� `�E/#z�)x� S232��� 1i� L�TEk@ PENDA�341 1D�3<*? �Mainten�ance Con%s B�? F"O,DNo UseM JOOnO�O�O�O�O2��2NPO;/" 1�9%�1CH=� 9�-Q		9Q_?!UD1:___�RSMAVAIL�/�/%�A!SR  �+��H�_�P�1�TVAL.&����P(.�YVL�}� �2i�� D��P 	�/_oUQ No�orci�o�g�o�o �o�o�o*,> tb������ ���:�(�^�L��� p�������܏ʏ �� $��H�6�X�~�l��� ��Ɵ���؟����� D�2�h�V���z����� ���ԯ
���.��R� @�b�d�v�����п�� �����(�N�<�r��i�$SAF_D?O_PULS. j0Qp����CA� ��/%�&0SCR �3�`4�X�
�0�0
	14�1IAIE���b vo$�6� H�Z�l�~�ߢߴ��߰�������HS"��2%���d1�(��8�rb��� @��"k�}���T�h� �J`���_ @��T7 �����#�~0�T D��0� Y�k�}����������� ����1CUg�y�O�Ef�p����  �5�;�o�� 1p��U�
�t���Di�������
  � ��*������ gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O7O<A���`OrO�O�O �O�O�O�O�O?O�_ ._@_R_d_v_�_�_�_�_�Q _�R0MJ To!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏJO��'�9�K� ]�o�������_ɟ۟ ����#�5�G�Y��_ �U�_�ҙ�����ϯ� ���)�;�M�_�m� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�;�?� q߮����������� ,�>�P�b�t�������������������Y��	�1234567�81h!B�!����F��� ��������������  ��;M_q ������� %7I[l*� ������// 1/C/U/g/y/�/�/�/ n��/�/	??-??? Q?c?u?�?�?�?�?�? �?�?O�/)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_O_ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �op_�o�o�o/ ASew���� �����o+�=�O� a�s���������͏ߏ ���'�9�K�]�� ��������ɟ۟��� �#�5�G�Y�k�}����������s�կ��w���0�L�CH�  Bpw�   ��=�2�� �} =�
~���  	�o�@ί��ǿٿ���r������@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖ�%� ����������&�8� J�\�n��������������"�Q�*�(����;�<M���D�~��  �]��w�*�Z򛱛�t C d�����*�`*���$SCR_GR�P 14*P�43� � }�*� 6��	 �
��<�+�*�'UC|@�Y�y�yD� W��!�y�	M-�10iA/7L �12345678k90��� 8���MT� � �
��	L��	Č� N
���Y���Dy�
M_	P������ ,���H�
 � ��1/@A/g/y/H���!T/�/P/�/3��+\���/B�S��,?�*2C4&Ad�R?  a@s�j5N?�7?��7�&2R��?}:&F@ F�`�2�?�/�? �?OO-OSO>OwObO �O=j1�2�O�O�O�O�DB��O�O;_&___ J_�_n_�_�_�_�_�_ o�_%o�5j�eSgxo6���uo�o�b�1�B�|3�oh0�4j96j9B� w�$0Y̯@HtA�Nhcu$�/�%pp�drsqA ����z�q�x�� �� (&� *�2�D�V�oz�e��������ECLVL ; ����iqp�Q@��L_DEF�AULT ���s�փH�OTSTR�qq���MIPOWER�F��H���WF�DO� �RVENT 1Ɂ�Ɂ� L!D?UM_EIP������j!AF_I�NE‧���!FIT}�֞����!-/�� ��F�!�RPC_MAIN�G�)��5���Y�VI�Sb�t����ޯ!�TPѠPUկ��d�ͯ*�!
PMON?_PROXY+���Ae�v��D���fe��¿!RDM_S�RVÿ��g���!#R,*ϑ�h��Z�K!
[�M����iI����!RLSYN�C����8����!�ROS|���4���>�!
CE�MOTCOM?ߓ�k-����!	S�CONSd�ߒ�ly���!SҟWASRCݿ��m���"�!S�USB�#n�n�!S#TMC��o]�� ���ѳ����,����P�V�ICE_KL� ?%d� (%�SVCPRG1S�����2�������oD����4������5D��6;@��7c h�����9����%������� ��0����X��� ��-���U���} ��� /���H/�� �p/���/��F�/ ��n�/��?�� 8?���`?��/�?�� 6/�?��^/�?��/X� j��q���#OhO��lO �O{O�O�O�O�O�O�O  _2__V_A_z_e_�_ �_�_�_�_�_�_oo @o+odoOo�o�o�o�o �o�o�o�o*< `K�o���� ���&��J�5�n� Y���}���ȏ���^�_DEV d���MC:�4����GRP �2d�
@�bx� 	� 
 ,V�ȡ�s�Z����� �������ߟ�� @�'�9�v�]�������@Я����۫Y��
@�ܯI�1�4�]��� j�����˿F�Ŀ�� %�7��[�B��f�x� ���!���A����ۿ D�+�h�Oߌ�s߅��� ������
���@�'�d�v��	y��^��� ��������%��I�0� Y��f�����8����� ������3��T7]�e�����)� �
�.@�dK �o��!�9���!/G/���R/ �/�/�/�/�/"�/�/ ??C?*?<?y?`?�? ��?�?�?�?�?�?-O OQO8OaO�OnO�O�O �O�O�O_�O)_;_"_ __�?�_�_L_�_�_�_ �_�_o�_7oo0omo To�oxo�o�o�o�o�o !x_E�oU{b �������� /��S�:�w�^�p������я�d �XƿZI6 r���@Z��0�+�A����d�BjBA�=��������B����AZ.�A����+�A.��Q�B�����5\��i6�A��u��'��ǎ%�Ꮛ�%�PEGA_BAR�RA_ESTEI�RA����X�T����?=��=�X��7
�?��>�A����?������&����������AxP��f���U�'A�j���´�B��:�<�3�����jB]+a��T��%�T�腯d�ʐ���>�p�c?��7�Գ�T@6��A�_���0n�����·�Ak���۸I�K9�FA�G�����B!v,�-���C3�����pBM�>�#�b��(�Y�������HX��?L!���Q��B���AJߤ�Xk�@f�D3��O�A���������Yw���.B��B�;��C�H�z�B�?���6���-Ϙ������n��=]����V@����?,����Ö� վ���eAk�������OY�A��ㇾ��AB��J�;%�C$�4�aƿBXZ�9���
���ߘ��~��� �ԭ(��?^_��-\¯ԡ���گ���+������������ߔ�mᢧ��*נ�6�C>�ԯb���z���
��BM����s��x�U<~�߯7@6|=��C��$�6��� N�@���b�G���L��}������x7���~K@����V�+A>r�rF���������Y@+�@��<B��|�A��F����B)���,o�?ɇ���~0��0~�6�Z� Q������������Aߍ�]ܖ�A����ܺ����2[�����>�ȥA���=�³�NB ��$�w?�d�j��to�7\��
�.�%��Z�����A������*�@Ve��B� ������YN�#���BD�	����9A����gB#
q��3��C4#���,?[BVM����COLO�CA_PRENS�����&//J/ 8/n/\/~/�/�/ �/�/�/ ??D?2?T? �/�/�?�/z?�?�?�? �?O
O@O�?gO�?0O �O,O�O�O�O�O�O_ ZO?_~O_r_`_�_�_ �_�_�_�_2_oV_�_ Jo8ono\o�o�o�o�o 
o�o.o�o"F4 jX��o��~� z���B�0�f�� ���V�����Џҏ� ��>���e���.��� ������̟Ο���X� =�|��p�^������� ��ȯ�D��T��H� 6�l�Z���~�����ۿ ���Ϡ��D�2�h� Vό�ο���|����� 
����@�.�dߦϋ� ��T߾߬�������� �<�~�c��,��� ��������D�)�;� �����\��������� ���@���4"D FX�|���� ��0@BT ����z��/ �,//</���/� b/�/�/�/�/?�/(? j/O?�/?�??�?�? �?�?�? OB?'Of?�? ZOHO~OlO�O�O�O�O O�O>O�O2_ _V_D_ z_h_�_�_�O�__�_ 
o�_.ooRo@ovo�_ �o�ofo�obo�o�o *N�ou�o>� ������&�h M�����n������� ��ȏ��@�%�d��X� F�|�j��������,� ��<�֟0��T�B�x� f���ޟï������� �,��P�>�t����� گd�ο�����(� �Lώ�sϲ�<Ϧϔ� �ϸ�������$�f�K� ���~�lߢߐ��ߴ� ��,��#�������D� z�h��������(� ���
�,�.�@�v�d� ������ ������� (*<r����� b����$ z�q�J��� ���/R7/v / j/�z/�/�/�/�/�/ */?N/�/B?0?f?T? v?�?�?�??�?&?�? OO>O,ObOPOrO�O �?�O�?�O�O�O__ :_(_^_�O�_�_N_p_ J_�_�_�_o o6ox_ ]o�_&o�o~o�o�o�o �o�oPo5to�oh V�z����( �L�@�.�d�R��� v������$���� �<�*�`�N���Ə�� �t�ޟp����8� &�\�����L����� گȯ����4�v�[� ��$���|�����ֿĿ ��N�3�r���f�T� ��xϮϜ������� ���Ͼ�,�b�P߆�t� ������ߚ����� �(�^�L���ߩ��� r����� �����$� Z������J������� ������b���Y�� 2�z����� :^�R�b� v����6� *//N/</^/�/r/�/ ��//�/?�/&?? J?8?Z?�?�/�?�/p? �?�?�?�?"OOFO�? mOO6OXO2O�O�O�O �O�O_`OE_�O_x_ f_�_�_�_�_�_�_8_ o\_�_Po>otobo�o �o�o�oo�o4o�o( L:p^��o�o �� ��$��H� 6�l�����\�ƏX� ֏��� ��D���k� ��4�������ҟ�� ��^�C����v�d� ��������ί��6�� Z��N�<�r�`����� �����󿪿̿��� J�8�n�\ϒ�Կ���� �����������F�4� j߬ϑ���Z��߲��� �������B��i�� 2������������ J�p�A����t�b��� ��������"�F��� :��Jp^��� ���� 6$ FlZ����� ��/�2/ /B/h/ ��/�X/�/�/�/�/ 
?�/.?p/U?g??@? ?�?�?�?�?�?OH? -Ol?�?`ONOpOrO�O �O�O�O O_DO�O8_ &_\_J_l_n_�_�_�O �__�_o�_4o"oXo Foho�_�_�o�_�o�o �o�o0T�o{ �oD�@���� �,�nS�����t� ��������Ώ�F�+� j��^�L���p����� ��ܟ��B�̟6�$� Z�H�~�l����ɯۯ ��������2� �V�D��z��������$�SERV_MAI�L  �����ʴOUTPUT�ո�@�ʴRV 2j� � � (r�������=�ʴSAV�E���TOP10� 2� d 6 rƱ���� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t������n�YPY��F�ZN_CFG f��=���J���GRP 2���g� ,B  � A �D;� �B �  B4~=�RB21I�oHELL��f�e�)�*�=�����%RSR��� ���&J5 G�k�������.�  ���/>/P/"\/ b�X/z"{ �U'
&"2�dh,g-�"E�HK 1S �/�/�/�/#?L?G? Y?k?�?�?�?�?�?�?��?�?$OO1OCO?OMM S�OD�FTOV_ENB�մ�e��"OW_R�EG_UI�O�IMIOFWDL~@��N�BWAIT��B�)��V��F��YTIM�E���G_VA԰_�A_�UNIT�C~Ve�L]C�@TRY�Ge��ʰMON_AL�IAS ?e�I%�he��oo&o8o Fj�_io{o�o�oJo�o �o�o�o�o/AS ew"����� ���+�=��N�s� ������T�͏ߏ�� ���9�K�]�o���,� ����ɟ۟ퟘ��#� 5�G��k�}������� ^�ׯ�����ʯC� U�g�y���6�����ӿ 忐����-�?�Q��� uχϙϫϽ�h����� ��)���M�_�q߃� ��@߹������ߚ�� %�7�I�[����� ����r������!�3� ��W�i�{���8����� ��������/AS e�����| �+=�as ��B����/ �'/9/K/]/o//�/ �/�/�/�/�/�/?#? 5?�/F?k?}?�?�?L? �?�?�?�?O�?1OCO UOgOyO$O�O�O�O�O �O�O	__-_?_�Oc_ u_�_�_�_V_�_�_�_�ooc�$SMO�N_DEFPRO�G &����Aa &�*SYSTEM*�obg $JO�0dRECALL �?}Ai ( ��}tpconn� 0 >10.1�09.3.23:�21152 2 �.*=�h1:11692 �a�`�a�o��o�o	v}7cop�y frs:or�derfil.d�at virt:�\tmpback�\�i�e�ofx~.�rmdb:*.*�2�oM���t2�xt:\�'��2A �a�s���q3�a%�7�I�R����� ,�P�a�s���� 3��N�ߟ����� ��L�]�o�����%�7� ʏۯ����$���H� 	�k�}�����=�ƟX� ���� ���D�ֿg� yό���/�¯T����� ���.�����c�u߇� ��5߾�P������� �ϸ�N�_�q���'� 9���������&߯� J�[�m���ߤ�?��� �������"��F��� i{���1��V� ���0���ew 
��7��R��/ ���a/s/�/��)/;/��/�/?>��:pickup�_barra_e�steira.tp�emp��!\?�n?�?<?/0torno9?��?�?�?z5�6lace�?��?�b�?dOvO�O};>�5sumir�?6O�J�O�O�O�?$D,3prens8?�O�Ok_ }_"71_C_K'Z_�_��_�Y=�Kfurad/_�_U?eowo
o�6��Csem_recep�@8oJo�o�o�oo#6co�o�o�oc�u� }:�5dr�op�bdefei�t�OIX��;8�z�t_1�I_�h�z���_23�E�W�0�������_3��ŏ ׏h�z��_1D�U� ��������ӟd��v����$SNPX�_ASG 2��������  01%����Я  ?���PARAM ��{�� �	���PӤ0Ө$�������OFT_�KB_CFG  �ӣ����OPIN_SIM  ���}����������RVNORDY_�DO  )�U����QSTP_DS�Bi��ϐ�SR� �� � �&#�D�O�O�:�T�OP_ON_ER�Rʿ��o�PTN �������A��RING_P�RMy�ܲVCNT?_GP 2��!���x 	����0`��#��Gߔ�VD���RP 1��"� 8Ѩ�*߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�}�z� ��������������
 C@Rdv�� ����	* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?[?X?j? |?�?�?�?�?�?�?�? !OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Losopo�o�o�o�o�o �o�o 96HZ l~��������� �2�D�V�`�P�RG_COUNT�J���{�ENBķ�}�M��L���_U�PD 1'�T  
k������"� K�F�X�j��������� ۟֟���#��0�B� k�f�x���������ү ������C�>�P�b� ��������ӿο�� ��(�:�c�^�pς� �Ϧϸ������� �� ;�6�H�Z߃�~ߐߢ� ���������� �2� [�V�h�z������ ������
�3�.�@�R� {�v������������� *SN`r���t�_INF�O 1�9Ҁ� 	 ���3��)X@�>��L9� C w�Bb?�	�;ӛ8�����,,MA�@��>>�` Ao�B @{w ?��� >�@���a ģ��C�Tp��1V�C3����"���3�����Y?SDEBUG����dՉ�SP_PwASS��B?+�LOG �.��  � a��  �с�U�D1:\;$�<"_MPCA-셽/�/��x!�/ 쁝&SAV D)��%d!l|"�%�(SV�+�TEM_TIME� 1D'�� 0�ν��
�',5�M7MEMBK  �сd d/�?��?�<X|Ҁ�3 @�?C�O:O�JLOmOzI�J�%@p1�O�O�O�O"3� __$_6_H_Z_l_ �n_�_�_�_�_�_�_�_o"o\�e1oVoho zo�o�o�o�o�o�o�o 
.@Rdv���O5SK�0�8��`�?���F.� e|�H2OJ�AJ�  @�C�A\O����(�O"�Oяb������p�O�"0� 	� ��0p�Z�l�~� r_���9�Ο������$�C�7og�y� ��������ӯ���	� �-�?�Q�c�u�����������T1SVG�UNSPD%% '�%��2MOD�E_LIM �a9"ܴ2�	� �D-۵ASK_OP�TION �9!�F�_DI ENB�  �5%f�BC�2_GRP 2!��u#o2��XB��C����ԼBCCFG 3#��*< #6���`�@I�4�Y� �jߣߎ��߲����� ����E�0�i�T�� x������������/��S�>�w����� t���u�����c��� 	B-f�.��4[  �������  02Dzh�� �����/
/@/ ./d/R/�/v/�/�/�/ �/�(���/?&?8?J? �/n?\?~?�?�?�?�? �?�?O�?4O"OXOFO hOjO|O�O�O�O�O�O �O__._T_B_x_f_ �_�_�_�_�_�_�_o o>o�/Voho�o�o�o (o�o�o�o�o(: Lp^���� ���� �6�$�Z� H�~�l�������؏Ə ��� ��0�2�D�z� h���To��ȟ���
� ��.��>�d�R����� ��z�Я������� (�*�<�r�`������� ��޿̿���8�&� \�Jπ�nϐϒϤ��� ���ϴ��(�F�X�j� �ώ�|ߞ��߲����� ���0��T�B�x�f� ������������� �>�,�N�t�b����� ������������: (^�v���� H���$HZ l:�~���� ���2/ /V/D/z/ h/�/�/�/�/�/�/�/ ?
?@?.?P?R?d?�? �?�?t�?�?OO*O �?NO<O^O�OrO�O�O �O�O�O�O__8_&_ H_J_\_�_�_�_�_�_ �_�_�_o4o"oXoFo |ojo�o�o�o�o�o�o �o�?6Hfx� �������v�&��$TBCSG_GRP 2$�u��  ��&� 
 ?�  Q�c�M���q��� �����ˏ��*�1��&8�d, ��F�?&�	 HCA;����b��?CS�B�I���<��V�>��ͪ�n��Ќ�ԝB��33Y3��Blt�������AÐ�fff�:��.�C����l�?����G�w�R���A&��̧�����@��I��-���
� X�u�@�R�����̻������	V3.0}0I�	mt7����*� �%��ֶY���@ff&� &�H�� N� �O�w  ����� �X�Ϙ�*�J21�'8���Ϥ�CFG -)�uB� E���+���d���#��#�I�W��pW� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ��������I�cp "4��gRw�� ����	-? �cN�r��&� �����/</*/ `/N/�/r/�/�/�/�/ �/?�/&??J?8?Z? \?n?�?�?�?�?�?�? O�? OFO4OjOXO�O �O`�O�OtO�O_�O 0__T_B_x_f_�_�_ �_�_�_�_�_�_,oo Poboto�o@o�o�o�o �o�o�o�o(L: p^������ �� �6�$�F�H�Z� ��~�����؏Ə��� �2��OJ�\�n���� ����������
� @�R�d�v�4������� ��ί����ү(�N� <�r�`���������ʿ ̿޿��8�&�\�J� ��nϐ϶Ϥ������� ��"��2�4�F�|�j� �ߎ����߀��� �� ��B�0�f�T��x�� �����������>� ,�b�P���������v� ������:(^ L�p�����  �$H6lZ |������/ �/ /2/h/�߀/�/ �/N/�/�/�/
?�/.? ?R?@?v?�?�?�?j? �?�?�?�?O*O<ONO OO�OrO�O�O�O�O �O�O _&__J_8_n_ \_�_�_�_�_�_�_�_ o�_4o"oXoFoho�o |o�o�o�o�o�o�/ $6�/�oxf�� ������,�>� ��t�b�������Ώ ��򏬏��&�(�:� p�^���������ܟʟ �� �6�$�Z�H�~� l�������دƯ���  ��D�2�T�z�h��� Jȿڿ������
� @�.�d�Rψ�vϬϾ� ���Ϡ������*� `�r߄ߖ�Pߺߨ��� �������&�\�J� ��n���������� ��"��F�4�j�X�z� |������������� 0B�Zl~(� ������, Pbt�D���8���   #� &0/"�$�TBJOP_GR�P 2*���  ?��&	H"O#,V,����� �z� =k%  Ȫ �� �� �$ �@ g"	 �C�A��&��SC���_%g!�"G���"k��/�+=��CS�?���?�&0%0CR  B4�'??J7��/�/?333�2Yx&0}?�:;��v 2R�1�0-1*20�6?��?20��7C�  �D�!�,� BL���OK:�Z�B_l  @pB@�� /s33C�1 �?gOO  A�zG�2jG��&)A)E�O�J;�}�|A?�ff@U@�1C�Z0zjO�Oz@ǰ��U�O�$ff�f0R)_;^;xCsQ?ٶ4)@�O�_tF��X_J\EU�_�V:�t-�Q(B�*@�Oo h�&-h$oZGLo6oDo ro�o~o8o�o�o�o�o 3�oRlVd(��V4�&`�q�%	V3.00m#Omt7A@�s*��l$!�'� E���qE���E��]\E�HF�P=F�{F�*HfF@D�F�W�3Fp?F��MF���F��MF��F��şF��F��=F���G�G.8��CW�RD3l)�D��E"���Ex�
E���E�,)FdR�FBFHFn� �F��F��M�F�ɽF�,
�GlGg!�G)�G=���GS5�GiĈ�;��
;�o��|& : @Xz�&/��&"�?��0�&=;-ESTP?ARS  (a �E#HRw�ABLEw 1-V) @�#R�7� � �R��R�R�'#!R�	�R�
R�R���!�R�R�R���RDI��`!��ԟ���
�r�Oz����� ����̯ޮ��Sx�^# <�����ÿտ��� ��/�A�S�e�wω� �ϭϿ�������;-w� {�_"��6��1�C�U� ��%�7�I�[���ҿNUM  �U`!� $  ���m���_CFG �.���!@H IM?EBF_TT}���^#��G�VE10m�H�z]�G�R 1/��O 8�" 2�� �A�  ��� ��������� �2�D� V�h�z����������� ��/
e@Rh v������� *<N`r� �����'/// ]/8/J/`/n/�/�/�/H�/r���_��t�@~��t�MI_CHA�NS� ~� !3DB/GLVLS�~�s��$0ETHERADW ?��w0�"���/�/�?�?l�$0R�OUTq�!�!��4�?�<SNMA�SKl8~�}1255.2E�s0OBOTO�s�t�OOLOFS_�DI}��%V9OR�QCTRL 0���#��MT�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo&l��OIo8omoq�PE_�DETAIJ8�JP�GL_CONFI�G 6�ᄀ�/cell/$�CID$/grp1qo�o�o/���?Zl~��� C���� �2�� V�h�z�������?�Q� ���
��.�@�Ϗd� v���������M���� ��*�<�˟ݟr��� ������̯@�}a�� �&�8�J�\���^o��c��`���˿ݿ�� �Z�7�I�[�m�ϑ�  ϵ����������!� ��E�W�i�{ߍߟ�.� �����������A� S�e�w����<��� ������+���O�a� s�������8������� '9��]o� ���F��� #5�Yk}������`�Us�er View ��i}}1234567890�//�,/>/P/X$� �cx/���2�U�/�/�/@�/??s/�/�3�/ b?t?�?�?�?�??�?�.4Q?O(O:OLO^OpO�?�O�.5O�O�O��O __$_�OE_�.6 �O~_�_�_�_�_�_7_�_�.7m_2oDoVoho zo�o�_�o�.8!o�o �o
.@�oagr� lCamera��o�� ��� �ޢE�*� <�N��h�z��������I  �v�)�� $�6�H�Z�l������ ����؟���� �2�Y��vP9ɟ~����� ��Ưد���� �k� D�V�h�z�����E�W� I5����� �2�D� �h�zό�׿������ ����
߱�W�ދ��X� j�|ߎߠ߲�Y����� ��E��0�B�T�f�x� ߁ulY��������� 
����@�R�d���� ������������W� i y�.@Rdv�/� ����* <N��W��i��� �����/*/</ �`/r/�/�/�/�/as9F/�/??1?C? U?�f?�?�?D/�?�?@�?�?	OO-O�j	�u0�?hOzO�O�O�O�O i?�O�O
_�?._@_R_ d_v_�_/OAO�p�{,_ �_�_oo)o;o�O_o qo�o�_�o�o�o�o�o �_�u���oM_q ���No���: �%�7�I�[�m�NE a����ˏݏ��� �7�I�[�������� ��ǟٟ����ͻp�%� 7�I�[�m��&����� ǯ�����!�3�E� 쟒�9�ܯ������ǿ ٿ뿒��!�3�~�W� i�{ύϟϱ�X����� H����!�3�E�W��� {ߍߟ�����������x����  �� L�^�p������������ ��    "�*�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/܄/�  
��( � �@�( 	 �/�/�/�/�/? ? 6?$?F?H?Z?�?~?�?�?�?�*2� � l�O/OAO��eOwO�O �O�O�O��O�O�O_ TO1_C_U_g_y_�_�O �_�_�__�_	oo-o ?oQo�_uo�o�o�_�o �o�o�o^opoM _q�o����� �6�%�7�~[�m� ��������ُ��� D�!�3�E�W�i�{� ԏ��ß՟����� /�A�S���w������ ��ѯ�����`�=� O�a�����������Ϳ ߿&�8��'�9π�]� oρϓϥϷ������� ��F�#�5�G�Y�k�}� �ϡ߳��������� �1�C�ߜ�y��� ����������	��b� ?�Q�c���������� ����(�)p�M�_q������0@� �������� ��#frh�:\tpgl\r�obots\m1�0ia4_7l.xml�Xj|��������.��/1/C/U/g/y/�/ �/�/�/�/�/�//? -???Q?c?u?�?�?�? �?�?�?�?
?O)O;O MO_OqO�O�O�O�O�O �O�OO _%_7_I_[_ m__�_�_�_�_�_�_ _�_!o3oEoWoio{o �o�o�o�o�o�o�_�o /ASew�� �����o��+� =�O�a�s����������͏ߏ�I ��<<  ?��4��,� N�|�b�������ʟ� Ο���0��8�f�L��~���������������(�$TPGL�_OUTPUT s9����� $�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ�@�ϳ�����$�����2345678901��� �2�D�V� ^����υߗߩ߻��� ��w����'�9�K�]���}g�������� o����1�C�U�g� ��u�����������}� ��-?Qc�� ������� );M_q	� ������%/7/ I/[/m///�/�/�/ �/�/�/�/?3?E?W? i?{??%?�?�?�?�? �?O�?OAOSOeOwO �O!O�O�O�O�O�O_��O� $$ Ӣ��OW=_o_a_�_�_ �_�_�_�_�_�_#oo Go9oko]o�o�o�o�o �o�o�o�oC5g}���������}@��"��? ( 	 iW� E�{�i�����Ï��ӏ Տ���A�/�e�S� ��w��������џ� ��+��;�=�O���s�����Ƹ  <<\ޯ�)�ͯ� )��M�_���ʯ���� <���ؿ��Ŀ� �~� $�V��BόϞ�x��� ��2ϼ�
ߤ���@�R� ,�v߈���p߾���j� ������<�߬�r� ���������� `�&�8���$�n�H�Z� �������������" 4Xj��R�� L����| Tf ��v�� 0B//�&/P/*/ </�/�/��/�/h/�/ ??�/:?L?�/4?�? ?n?�?�?�?�? O^? �?6OHO�?lO~OXO�O �OO$O�O�O�O_2_ __h_z_�O�_�_J_��_�_�_�_o.o��)�WGL1.XM�L�cm�$TPOFF_LIM Š|�p���qf�N_SVy`  ��t�jP_MON7 :���d�p��p2miSTRT?CHK ;���f�~tbVTCOM�PAT�h*q�fVW�VAR <�m\Mx�d  e��p�bua_DE�FPROG %��i%COLO�CA_MESA_?IRVISI�`~�rISPLAY�`��n�rINST_M�SK  �| ~�zINUSER ��tLCK)��{QUICKME�pO��roSCREl���~+rtpsc�t�)������b��_��S�Tz�iRACE_�CFG =�i�Mt�`	nt
?�~�HNL 2>�z���T{ zr@�R�d��v���������К�I�TEM 2?,�� �%$1234?567890�%�  =<�C�U�]��  !c�k�wp '���ns�ѯ5���� k������j�ů��� ����A�1�C�U�o�y� 󿝿I�oρ�忥�	� �-ϧ�Q���#�5ߙ� A߽�����e߳���� ��M���q߃�L��g� �ߋ����%�w� � [���+�Q�c���o� �������3��� {�;������G_�� ��/�Se.� I�m�� �=�a/3/�� ����k//�/�/ �/]/?�/�/�/?�/ u?�?�??�?5?G?Y? �?+O�?OOaO�?mO�? �?�OO�OCO__yO +_�O�Ox_�O�_�O�_ �_�_?_�_c_u_�_o �_Wo}o�o�_�oo)o ;o�o�oqo1C�oO �o�o��%��@[��Z��S��@��_��  �ے_� ����y
� Ï�Џ����UD1:\����q�R_GRP 1�A �� 	 @�pe�w�a���������ߟ͞�����ّ�>�)�b�M�?�  }���y�����ӯ ������	��Q�?� u�c���������Ϳ��	-���o�SC�B 2B{�  h�e�wωϛϭϿ��������e�UTORIAL C{��@��j�V_CONFIG D{����������O�OUTPUT� E{�����������%�7�I� [�m�������� ������%�7�I�[� m�������������� ��!3EWi{ �������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/��/??'?9?K? ]?o?�?�?�?�?�?�/ �?�?O#O5OGOYOkO }O�O�O�O�O�O�?�O __1_C_U_g_y_�_ �_�_�_�_�O�_	oo -o?oQocouo�o�o�o �o�o�_�o); M_q����� �yߋ����-�?�Q� c�u���������Ϗ� ��o�)�;�M�_�q� ��������˟ݟ� � �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i�{������� ÿտ���
��/�A� S�e�wωϛϭϿ��� ������+�=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� �����������1 CUgy���� ���	-?Q cu��������/�x��� $/6/ !/a/��/�/ �/�/�/�/�/??'? 9?K?]?�?�?�?�? �?�?�?�?O#O5OGO YOkO|?�O�O�O�O�O �O�O__1_C_U_g_ xO�_�_�_�_�_�_�_ 	oo-o?oQocot_�o �o�o�o�o�o�o );M_q�o�� ������%�7� I�[�m�~������Ǐ ُ����!�3�E�W� i�z�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'��9�K�]�o�~��$T�X_SCREEN� 1F8%  �}�~���������
����m&�� \�n߀ߒߤ߶�-�?� �����"�4�F��j� �ߎ���������_� ���0�B�T�f�x��� ���������� ��>��bt��� �3�W(: L^������ ��e/�6/H/Z/�l/~/�//�/�$U�ALRM_MSG� ?�����  �/���/�/)??M?@? q?d?v?�?�?�?�?�?��?O�%SEV  ��-EF�"EC�FG H����  ��@� � AuA   B���
 O���ŨO �O�O�O�O__&_8_�J_\_jWQAGRP �2I[K 0��	� �O�_� I_B�BL_NOTE �J[JT�G�l������g@~�RDEFPRO� �%�+ (%C�OLOCA_ME�SA_IRVISION�_%OVoAo zoeo�o�o�o�o�o�o��o@�[FKE�YDATA 1K<�ɞPp jG���_������z�,(����([ INST ]'�)�v@CROS�}�d�?REL  T��� CHOICEB����[EDCMD Ə��&��J�1�n� ��g�����ȟڟ������"�4��X��z���/frh/gu�i/whitehome.pngd�`����Ưدꯀ{�inst���/�A��S�e���  |�pgmacro������ȿڿ�{�gkarel��(�:�L�^�p���clos��ϯϠ����������{�edcmd�3�E��W�i�{���{�arwrg��������� �߁��)�;�M�_�q� ������������ ��%�7�I�[�m��� �������������� 3EWi{�� �����/A Sew��r��� ���/!/(E/W/ i/{/�/�/./�/�/�/ �/??�//?S?e?w? �?�?�?<?�?�?�?O O+O�?OOaOsO�O�O �O8O�O�O�O__'_ 9_�O]_o_�_�_�_�_ F_�_�_�_o#o5o�_ Goko}o�o�o�o�oTo �o�o1C�og y����P�� 	��-�?�Q��u����������Ϗj�܋�u�܏�(�s���Q�c�r�,I���A�O?INT  ]����? OOK Tß�~}�NDIRECܟ��  CHOIC�E�����UCHUPG�H�s���~����� ߯�د���9�K�2� o�V�������ɿ���whitehom ����%�7�I�X���poin�ߍϟϱ������d�i/look��#�5�G�Y����i/indirec|Ϙߪ߼�����g�choic���� ��2�D�V�h�k�touchup�ߠ���������g�arwrg ��"�4�F�X�j�a��� ����������w� 0BTfx�� �����,> Pbt���� ��/�(/:/L/^/ p/�//�/�/�/�/�/  ?׿�/6?H?Z?l?~? �?�/�?�?�?�?�?O �?2ODOVOhOzO�O�O -O�O�O�O�O
__�O @_R_d_v_�_�_)_�_ �_�_�_oo*o�_No `oro�o�o�o7o�o�o �o&�oJ\n ����E��� �"�4��X�j�|��� ����A�֏����� 0�B�яf�x������� ��O������,�>��<L������u�����q���ͯ��,������"�	� F�X�?�|�c������� ֿ������0��T� f�Mϊ�qϮϕ����� �����,�>�?b�t� �ߘߪ߼�˟����� �(�:�L���p��� �����Y��� ��$� 6�H���l�~������� ����g��� 2D V��z����� c�
.@Rd �������q //*/</N/`/��/ �/�/�/�/�/�//? &?8?J?\?n?�/�?�? �?�?�?�?{?O"O4O FOXOjO|OSߠO�O�O �O�O�OO_0_B_T_ f_x_�__�_�_�_�_ �_o�_,o>oPoboto �oo�o�o�o�o�o �o:L^p�� #���� ��� 6�H�Z�l�~�����1� Ə؏���� ���D� V�h�z�����-�ԟ ���
��.���R�d� v�������;�Я��� ��*���N�`�r���Ж������@���>�@������ 	��+�=��,)�n� !ߒ�y϶��ϯ����� �"�	�F�-�j�|�c� �߇����߽������ �B�T�;�x�_��� �O��������,�;� P�b�t���������K� ����(:��^ p����G��  $6H�l~ ����U��/  /2/D/�h/z/�/�/ �/�/�/c/�/
??.? @?R?�/v?�?�?�?�? �?_?�?OO*O<ONO `O�?�O�O�O�O�O�O mO__&_8_J_\_�O �_�_�_�_�_�_�_�� o"o4oFoXojoq_�o �o�o�o�o�o�o�o 0BTfx�� ������,�>� P�b�t��������Ώ ������(�:�L�^� p��������ʟܟ�  ����6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z����� -�¿Կ���
�ϫ� @�R�d�vψϚ�)Ͼπ��������*�`�,��`���U�g�y�Qߛ߭߇�,���ߑ����&�8� �\�C���y��� ���������4�F�-� j�Q���u��������� ���_BTfx �������� ,�Pbt�� �9���//(/ �L/^/p/�/�/�/�/ G/�/�/ ??$?6?�/ Z?l?~?�?�?�?C?�? �?�?O O2ODO�?hO zO�O�O�O�OQO�O�O 
__._@_�Od_v_�_ �_�_�_�___�_oo *o<oNo�_ro�o�o�o �o�o[o�o&8 J\3����� ��o��"�4�F�X� j��������ď֏� w���0�B�T�f��� ��������ҟ����� �,�>�P�b�t���� ����ί�򯁯�(� :�L�^�p�������� ʿܿ� Ϗ�$�6�H� Z�l�~�Ϣϴ����� ����ߝ�2�D�V�h� zߌ�߰��������� 
��.�@�R�d�v�ﴚ�qp���qp���������������,	N�r� Y������������� ��&J\C�g �������" 4X?|�m� ����/�0/B/ T/f/x/�/�/+/�/�/ �/�/??�/>?P?b? t?�?�?'?�?�?�?�? OO(O�?LO^OpO�O �O�O5O�O�O�O __ $_�OH_Z_l_~_�_�_ �_C_�_�_�_o o2o �_Vohozo�o�o�o?o �o�o�o
.@�o dv����M� ���*�<��`�r� ��������̏���� �&�8�J�Q�n����� ����ȟڟi����"� 4�F�X��|������� į֯e�����0�B� T�f�����������ҿ �s���,�>�P�b� �ϘϪϼ������� ���(�:�L�^�p��� �ߦ߸�������}�� $�6�H�Z�l�~��� ����������� �2� D�V�h�z�	��������������
�}�����5@GY1{�g,y �q���< #`rY�}�� ���/&//J/1/ n/U/�/�/�/�/�/�/ �/ݏ"?4?F?X?j?|? ���?�?�?�?�?�?O �?0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�_�_'_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o $�oHZl ~��1���� � ��D�V�h�z��� ����?�ԏ���
�� .���R�d�v������� ;�П�����*�<� ?`�r����������� ޯ���&�8�J�ٯ n���������ȿW�� ���"�4�F�տj�|� �Ϡϲ�����e���� �0�B�T���xߊߜ� ������a�����,� >�P�b��߆���� ����o���(�:�L� ^�������������� ��}�$6HZl ��������y  2DVhzQ��|�Q�����������,�/./�/R/9/v/ �/o/�/�/�/�/�/? �/*?<?#?`?G?�?�? }?�?�?�?�?OO�? 8OO\OnOM��O�O�O �O�O�O�_"_4_F_ X_j_|__�_�_�_�_ �_�_�_o0oBoTofo xoo�o�o�o�o�o�o �o,>Pbt� ������� (�:�L�^�p�����#� ��ʏ܏� ����6� H�Z�l�~������Ɵ ؟���� ���D�V� h�z�����-�¯ԯ� ��
����@�R�d�v� �������Oп���� �*�1�N�`�rτϖ� �Ϻ�I�������&� 8���\�n߀ߒߤ߶� E��������"�4�F� ��j�|������S� ������0�B���f� x�����������a��� ,>P��t� ����]� (:L^���� ���k //$/6/ H/Z/�~/�/�/�/�/h�/�/���+������?'?9=?[?m?G6,YO�?QO �?�?�?�?�?OO@O RO9OvO]O�O�O�O�O �O�O_�O*__N_5_ r_�_k_�_�_�_�_�� oo&o8oJo\ok/�o �o�o�o�o�o�o{o "4FXj�o�� ����w��0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� ����(�:�L�^�p� �������ʯܯ� � ��$�6�H�Z�l�~��� ���ƿؿ���ϝ� 2�D�V�h�zό�ϰ� ��������
���_@� R�d�v߈ߚߡϾ��� ������*��N�`� r����7������� ��&���J�\�n��� ������E������� "4��Xj|�� �A���0 B�fx���� O��//,/>/� b/t/�/�/�/�/�/]/ �/??(?:?L?�/p? �?�?�?�?�?Y?�? O�O$O6OHOZO�$U�I_INUSER  ���{A��  �[O_O_MENH�IST 1L{E�  (� �@��(/S�OFTPART/�GENLINK?�current=�menupage?,153,1�O_�_1_C_�'�O�N7�1�@BARRA_ESTEIRA�O��_�_�_�3)X_�Ee�dit�BMAIN>�PLACE0�_o .o@oK_�_�I2�Ao��o�o�o�o�Opo,148,2�o/A�S�9�o�^COL�OCA�@SA_I?RVISIOa�8����� i�o 	"�4�F�X����O`����ď֏�6���0 �A����"�4�F�X� j�m���������ȟڟ �{��"�4�F�X�j� ��������į֯�w� ��0�B�T�f�x�� ������ҿ������ ,�>�P�b�t�ϘϪ� ����������(�:� L�^�p߂߅�#߸��� ���� ���6�H�Z� l�~���������� ������D�V�h�z� ����-���������
 ��@Rdv�� );���* �N`r���� ���//&/8/� \/n/�/�/�/�/E/�/ �/�/?"?4?F?�/j? |?�?�?�?�?S?�?�? OO0OBO�?fOxO�O �O�O�O�OaO�O__ ,_>_P_;t_�_�_�_ �_�_�_�Ooo(o:o Lo^o�_�o�o�o�o�o �oko $6HZ l�o������ y� �2�D�V�h�� ������ԏ�������.�@�R�d�v�aX��$UI_PANE�DATA 1N�������  	�}  �frh/cgtp�/flexdev�.stm?_wi�dth=0&_h�eight=10�ԐŐice=TP�&_lines=�3Ԑcolumnws=4Ԑfonܐ�4&_page=/doubŐ1��\V?)  rim#�L�  ��c�u������� ��$�ϯ�گ���;� M�4�q�X�������˿������%�\V�� �   nP��]���ʟܝ�2����2/�-�ual����_��"�4� F�X�j�ώ�u߲��� ���������B�)� f�M������3�E�  ���� ���*�<�N�`��� ���Ϩ��������� i�&8\C�� y������ 4Xj=���� ������� /S $/��H/Z/l/~/�/�/ 	/�/�/�/�/�/ ?2? ?V?=?z?a?�?�?�? �?�?�?
O}�@ORO dOvO�O�O�?�O1/�O �O__*_<_N_�Or_ Y_�_}_�_�_�_�_�_ o&ooJo1ono�ogo �oO)O�o�o�o" 4�oXj�O��� ���O��0�B� )�f�M����������� ���ݏ��>��o�o ���������Ο��3� �w(�:�L�^�p��� 韦�����ܯï �� ��6��Z�A�~���w� ����ؿ�]�o� �2� D�V�h�z�Ϳ����� ������
��.ߕ�R� 9�v�]ߚ߬ߓ��߷� �����*��N�`�G�����	�������������"�)��G���6� s�����������4��� ����K2oV ���������#�����$UI�_POSTYPE�  �� 	 /�U�QUICKMEN  ds�W�RESTORE �1O� � ��� /#���m+/T/f/ x/�/�/?/�/�/�/�/ ?�/,?>?P?b?t?/ �?�?�??�?�?OO (O�?LO^OpO�O�O�O IO�O�O�O __�?_ 1_C_�O~_�_�_�_�_ i_�_�_o o2o�_Vo hozo�o�oI_So�o�o Ao�o.@Rd �����s�� �*�<��oI�[�m�� ����̏ޏ�����&� 8�J�\�n��������xȟڟ�SCRE��?�u1�sc�u2�3��4�5�6�7r�8��TAT`�� ��MUScER�����ks����3��4��5��6ʨ�7��8��UND�O_CFG P�d����UPDX�����Non�e���_INFOW 1Q�<��0%��W���E���i� ��������տ��� :�L�/�pς�eϦύ�)�OFFSET Td@���{�� ����	��-�Z�Q�c� �߇ߙ��ϝ�������  ��)�V�M�_�q��������
���t���)�WORK U4�����A�S������UFRAME � ���&�RTO?L_ABRT��$�μ�ENB����GR�P 1V��Cz  A��� +=Oas��ĸ��U������MS�K  �<���N6��%4��%��)���_EVN������>�2W��
 }h��UEV���!td:\ev�ent_user\-�C7���}�YF��SP���spotweld�!C6����!�Z/�/:' �H/~/l/�/�/�/�/ -?�/Q?�/? ?�?D? �?h?z?�?O�?)O�? �?OqO`O�O@ORO�O vO�O_�O�O7_�O[_h_Z]W+�2X��F��8V_�_�_ �_ �_o�_,o>ooboto Oo�o�o�o�o�o�o �o:L'p�]�����$VARS_CONFI��Y�� FP{����|CCRG�\P��>�{�t�D�� BH� pk�a�Ce�� ��}�?����C,&Q=��ͩ�Am �MR2b��'�	}�	��@��%1: SC130EF2 *�����{�����X� �e5}�����A@k�;C�F� w�Q�[���|���������D�T����\�ϟ� �\� B���;�e�@�ǟ`����� S�����̯���ۯ� &�}��\�G�Y���E����ȿ�TCC�c�
��������pG�F�pgd���-�23456789017�?��ׁ$���4�v�Nm�� ��϶�BW�����i�}�?:�o=LA�څ �6�@�6�ͿZ���i�7����(��W���-� ]�X�jĈߚߕϳϹ� ��������%�7�I� r�m�ߨ�ߵ����� �����8�3�E�W�� ����}����������� ��/�A�S�e�w���MODE��t ��RSLT e�|k�%"zς��;� 1��d��`��SELEC��c�}�	IA_WO�P�f �� >W,		�����>�G�P ������RTSYNCS�E� ��$�	#WINURL ?*ـ�;\/n/�/�/��/�/�uISION�TMOU���A# ���%�gSۣ��SۥP�� �FR:\�#\D�ATA\�/ �߀ MC6LO�G?   UD�16EX@?\�'� B@ ����2T1Gabri�el_Faria�k?P5�?�?������ n6  ����GV�2\� -�|�5��   ���Z�@U058TRACINj?��*B{Rd_C�p��D #A`{2��'$�"��h#� (�kI�Mw��O �O�O�O�O1__U_C_�]_g_y_�_�_�_�(SKTA� i��@���o0oI:$obo�%_kGE�j#��~@� �
�\��btgH�OMIN�kS����`�2,,���CWǖBveJMP�ERR 2l#�
  QoI:��"� 4Fwj|����������&%S-_g0RE�m�^۴�LEXdn�1�-ehoVMPHA�SE  �e׃�BޱOFF _E�NB  �$V�P2�$oSۯR��x�c C;�@ ��@�;���?s33'D*AA��]� �P�0ޱ�`r}�XC ��܅���\A-۟E ������#� 5�������������}� ���������c�X� ��A�����ϯ�+�� ߿��M�B�q���x� �Ϲ���Ϸ������� 7�I�;�m�b�)ߣ�E� �ߡ߳�����3��� W�L�{ߍ��ߑ��� �������/�$�6�e� W���c�y��������� �����O���?M _q������� '9�=7Is� �����/m�/%/3/E/s�TD__FILTE�`s�kg �x2�`��� �/�/�/�/�/	??-? ??Q?�6�/~?�?�?�?��?�?�?�?O OoiS�HIFTMENU� 1t}<5�% 5�~O)�\O�O�O�O�O �O�O�O'_�O_6_o_�F_X_�_|_�_�_�_�	LIVE/SN�AP�Svsflsiv���_�z`/ION ҀU
`bmenu&o+o�_�oP�oV"<E�uz��4IkMO�v���zq��WAITDINEND  �ec��b��fOKوOUT��hSDyTIM.du��o|G�} #�{C�zb�z�x�RELE��ڋxT�M�{�d��c_A�CT`و��x_D?ATA wz����%  EGA_B�ARRA_EST�EIRA�o6Ex�R�DIS
`E��$�XVR�ax�n��$ZABC_GRoP 1yz���� ,�2̏.MZ�D��CSCH�`zd���aP@�h@�IP�b{'����şן�[�MPCF__G 1|'���A0�r�8��� �}'���p�s� 	|(���  <l0�  ��  ����5�>�����?��5�`���?5�U������C�Tp���1V�>w�@3�>�?|�/�Q���6 `��@Q�>���`���� ��˯ݯ����o�p��w���� /��C3����"��3��˿ݸĸ� �	��1�?�i���'�9�0?�Q��	��`�~����_CYLI�ND~!� ��� ,(  * .�?ݧ+�h�Oߌ�s� ��������(�	� x�-��&�c�߇�� ������j�P����)���~�_�q��� �2�'��� �&���� ������&��I��cA���SPH�ERE 2��� �������A� T/A��e�� ����/N` =/�a/H/Z/�/��/��/�/�ZZ� � �f