��   g�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����BIN_CFG_�TX 	$EN�TRIES  �$Q0FP?N�G1F1O2F2�OPz ?CNET�G  �DHCP�_CTRL. � 0 7 ABL�E? $IPUS~�RETRAT��$SETHOS�T��NSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM�� !� FT�� @� LOG_�8	,CMO>$�DNLD_FIL�TER�SUBD�IRCAPC  �D��8 . 4� H{ADDR�TYP�H NG#TH���z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~�OMGDEV������PINFO~�  $�$$TI� �R�CM+T �A$( /�QSI�Z�!S� TAT�US_%$MAI�LSERV $�PLAN� <$�LIN<$CLyU��<$TO�oP$CC�&FR�&�YJEC|!Z%E�NB � ALA5R:!B�TP,�#�,V8 S��$VkAR�)M�ON�&����&APPL�&P�A� �%��'POR��Y#_�!�"ALE�RT�&i2URL �}Z3ATTA�C��0ERR_T7HROU3US�9H!��8� CH- c%�4M�AX?WS_|1;��1MOD��1AI�  �1o (�1�PWD  � LAط�0�ND�1TR=YFDELA-C�0<G'AERSI��1vQ'ROBICLK_HqM 0Q'� XML+ �3SGFRMU3T̑ !OUU3 G_�-COP1�F33�A�Q'C[2�%�B_AU��� 9 R�!UP=Db&PCOU{!�C�FO 2 
�$V*W�@c%AC�C_HYQSNA�U�MMY1oW2"$D�M*� $DI�S�� SM�	 l5�o!�"%Q7�IZP�%� �V�R�0�UP� _DL�VSPAR!#�PN,#
3 �_�R!�_WI�CTZ_I�NDE�3^`OFF,� ~URmiD�)c��   t 9Z!`MON��c�D��bHOUU#E�%A�f�a�f�a�fLOsCA� #$NS0oH_HE���@�I�/  d8`A�RPH&�_IPFF�W_* O�F``�QFAsD90�VHcO_� 5R42PSWq�?�TEL� �P���90W�ORAXQE� L�V�[R2�IC�E��p� �$cs G  �q��
���
�p�PS�A�w[# 0�	�Iz0�AL��' �
���F���P��!�p��i��$� 2Q������������ Q���!�q�����$� _FLTR � �\� ��
��������$Q��2��7rSH`D +1Q� P㏙�f���ş��韬�� П1���=��f���N� ��r�ӯ�������ޯ �Q��u�8���\��� ����󿶿�ڿ;��� _�"�XϕτϹ�|��� ��������6�[�� �Bߣ�f��ߊ��߮� ��!���E��i�,�� P�b���������� /���(�e�T���L���l��z _LUA1�_x!1.��0���p���1��p�25c5.0��r��n���2����d %7I[3e��� ����[4���T'9[5U��� {���[6���@D �//)/s��Q�ȁMA��M?A� ����� Q� ��u.<�/?&?�/J?\? n?A?�?�?m�P�?�? �?�?�?O.O@OROOvO�O�Ou.kOl�q���O�L
ZDT ?StatusZO�O�5_G_Y_n�}iR�Connect:� irc{T//alert^�_�_�_ �_mW#_oo,o>oPo�bot�^�d~2g���go�o�o�o�o�o�o 	-?Qcul��$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5_2e036�`(�_��_���"�p�1!W��(��"S��J�E�� X��C� ��,$ ���W���ˏ��� ֏��%��I�0�m�� f�����ǟ�������h!��u�R����n� DM_�!�����SMTP_CT�RL 	����%����DF���ۯt�@ʯ��'��Lz�N�B�!
j��y�q�u����Ԙ��#L��USTOM dj������  ����$TCPIPd��j��H�%�"�EL������!���H!�TP��j�rj3_tp�b;���~i�!KCLG��L�i���5�!CR�T�ϔ����"u�!�CONS��M��[�ib_smon����