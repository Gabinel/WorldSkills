��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@&8&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	�>&USRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  w0�aIRTs1�	o`'2 L1��L1��R�	 �,��?���a�1`�b�ba ���a�� ��  ����
 ��a�o�o1CU �oz�� ���c�
��.� @�R��v��������� Џ�q���*�<�N� `��������̟ޟ m���&�8�J�\�n� ��������ȯگ�{� �"�4�F�X�j����������Ŀֿ���`�TPTX��p���/�` s����$/soft�part/gen�link?hel�p=/md/tpmenu.dg�� �ϨϺ��υ����� &�8�J���n߀ߒߤ� ����W������"�4� F�X���|�����������a�f�oC ($p�-����T�?�x���a�a�� �c���c����l��cP�g�e�a�a�dh���a2�h�	f���%�������`����`  ���f eOp��h#h��F�bc Xc�B 1�)hR \� _�� ;REG VED]����wholem�od.htm�	s�ingl	do�ub tri�p8browsQ�����u ���//@/��|�dev.s�l�/3� 1�,	t �/_�/;/i/??/?��/S?e?w?�?�?�?� ��?�?OO%O�7OIO[OmOO�E @ �?�O�O�O�O�O_�F �	�?�?;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omooM'�o �o�o�o�o�o+ =Oas���� �����?>�P�b� t���������Ώ���O �����L�^�_'_ �������ş���� �6�1�C�U�~�y��� ��Ư��ӯ�o��� -�?�Q�c�u������� ��Ͽ����)�;� M�_�-��ϬϾ����� ����*�<�7�`�r� A�Sߨߺ�q���i�� ���!�J�E�W�i�� ������������"� �/���O�I�w����� ����������+ =Oas���� ���,>Pb t���߼��� //�����^/Y/k/ }/�/�/�/�/�/�/�/ ?6?1?C?U?~?y?�? Y��?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__�R_ d_v_�_�_�_�_�_�_ �_�o*o�_o`oro��j�$UI_TO�PMENU 1�K`�aR� 
d�a*Q)�*default�5_]*lev�el0 * [	 #�o�0�o�'rtpio[23�]�8tpst[1[x)w9�o	�=�h58E01_�l.png��6menu5�y�p�C13�z��z	�4���q��]������� ��̏ޏ)Rr���+��=�O�a���pri�m=�page,?1422,1h��� ��şן����1��C�U�g���|�class,5p������ɯۯ�����13���*�<�N�`�r���|�53������ҿ�����|�8��1�C� U�g�y����ϯ���������"Y�`�a�o/߀�m!ηq�Y��avt�yl}Tfqmf[0�nl�	��c[164[w��59[x�qG�Ly��tC8�|�29� �o�%�1���{��m� �!�����0�B��� f�x���������o���80��'9K~���2P���� �\��'9K ������������1��/$/6/H/�Z/U�|�ainedi'ߑ/�/�/�/�/�P�config�=single&>|�wintp���/ $?6?H?Z?	�ߐ??�>��gl[57�ٳ q��?�;gp�08�ݲ0A7I�?F��F2JO[6�:�?)O�O�x �6� �4s�x�O ���$��`�o�H_Z_ l_~_�_�_Q��_�_�_ �_o o�_DoVohozoЌo�o�o�!;�$dokub5o��13���&dual�i38���,4�o&�o9 �o�n�o�a8��� Ao����&�8��%�3L=}!��o�b8 @���������z����(�:��+:T��i48,2o��b{����ʟ {?�;�M�sc���;���s�� �}����e�u��X��@�F7L���`�O��2�h�z�6e�u7������Ͽ���̏�27��G�Y�k�}Ϗ�� 0�s���������!�1�M�_�q߃� ������������� ��7�I�[�m���� ����������!�����6(�]�o��������$��746������)�C�ߟT�	�TPTX[209�<Aw2IHJ���Bw1H�]H�����02��A#��[Ttv`��O�L#_�0� \��5S[��treeview�3v�3��~�381,26M/_/q/0� �/�/�/�/�/�/~/? %?7?I?[?m?�o/(���o5%���?�?�?�AD�?\1~��?8"2�� eOwO�?�?(}�LEK� �O�O_�O��8@�ONOa_s_�_��6_d�E_ �_�_�_oV�#_���_ �Sooo�o�oB�o�o ��oA�oq+ =Oas��o�� �����(�9��� Q�x���������ҏ? ����,�>�P�ߏt� ��������Ο]���� �(�:�L�^�ퟂ��� ����ʯܯk� ��$� 6�H�Z��l������� ƿؿ�y�� �2�D� V�h����Ϟϰ����� �ϕo�o��o@ߧE� c�u߇ߙ߽߬����� O����)�<�M�_�q� ���W��������� &�8���\�n������� ��E�������"4 ��Xj|���� S��0B� fx����O� �//,/>/P/�t/ �/�/�/�/�/]/�/? ?(?:?L?��߂?1� �?���?�?�?�?O $O5OGO�?SO}O�O�O �O�O�O�O�O��2_D_ V_h_z_�_�_�/�_�_ �_�_
oo�_@oRodo vo�o�o)o�o�o�o�o *�oN`r� ��7����� &��J�\�n������� ��E�ڏ����"�4� ÏX�j�|�������a? s?蟗?�sO_/�A� S�e�w���������� �����,�=�O�a� #_������ο��=� �(�:�L�^�pς�� �ϸ������� ߏ�$� 6�H�Z�l�~�ߐߴ� ����������2�D� V�h�z�������� ����
����@�R�d� v�����)����������ƚԔ*de�fault%��*level8��ٯw���? tpst[1]�	��y�tpioG[23���u����J\men�u7_l.png�_|13��5Ж{�y4�u6 ���//'/9/K/]/ ���/�/�/�/�/�/j/ �/?#?5?G?Y?k?�"�prim=|p�age,74,1�p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_ �_�_�__B6o9o�Ko]ooo�o`�$U�I_USERVI�EW 1֑֑�R 
����o��o�o[m �o'9K] � ����l��� #�5��oB�T�f���� ��ŏ׏鏌���1� C�U�g�
��������� ӟ~�����v�?�Q� c�u���*�����ϯ� 󯖯�)�;�M�_�
��*zoomr�?ZOOMIN�q� �ؿ���� �ÿD� V�h�zό�/ϰ����������Z*maxr�es��MAXRES��	ߧ�p߂ߔߦ� ��[����� ��$��� H�Z�l�~��;ߡ�� ��3���� �2�D�V� ��z���������e��� ��
.��;Q_ �������� *<N`�� ���w��/o 8/J/\/n/�/#/�/�/ �/�/�/�/?"?4?F? X?/i?w?�?�/�?�? �?�?OO�?BOTOfO xO�O-O�O�O�O�O�O �?__'_�Ob_t_�_ �_�_M_�_�_�_oo (o�_Lo^opo�o�o7a