��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� �G_~�0COUPLE, �  $�!PP�V1CES0�!H1��!�PR0�2	 �� $SOFT��T_IDBTO�TAL_EQ� �Q1]@NO`BU SP?I_INDE]uE�XBSCREENu_�4BSIG�0�O%KW@PK_�FI0	$T�HKY�GPANE�hD � DUMM�Y1d�D�!U4� Q!RG1R�
 � $TIT1d ��� 7Td7T� �7TP7T55V65V7*5V85V95W05W>W@�A7URWQ7UfW1pW1zW1�W1�W 6P~!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$Nb_OPT�2 � �ELLSETUP�  `�0HO��0 PRZ1%{cM�ACRO�bREP	R�hD0D+t@��bl{�eHM MN�yB
1�UTOB �U�0 �9DEVIC4ST	I�0�� P@13�r�`BQdf"VAL�#ISP_UNI��#p_DOv7IyFR_F�@K%D13�x;A�c�C_WA?t��a�zOFF_@N.�DEL�xLF0q8�A�qr?q�pF�C?�`�A�E�C#��s�ATB�t�d��MO� �sE �� [M�s��2�R;EV�BILF��1�XI� %�R � � OD}`j�_$NO`M� +��b�x�/�"u��� ����!X�@D�d p E R�D_Eb��$F�SSB�&W`KBD�_SE2uAG� G
�2 "_��B�� V�t:5`ׁQC �a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR�B�IGALLOW�� (KD2�2�@VAR5�d!�AB �e`BL[@S � !,KJqM�H`S�pZ@�M_O]z����CFd X�0G�R@��M�NF�LI���;@UIR�E�84�"� SWIYT=$/0_No`S�"�CFd0M� =�#PEED��!��%`���p3`J3tV�&$E�..p`L�>�ELBOF� ��m��m�p/0��CP�� F�B����1���r@1J1E_y_T>!Բ�`��g����G� �0WARNMxp�d�%`��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqM��� R�r$ORIأ.&ӧRT�SF\g CHGV0I�Ep�T��PA�I{��T�!��� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5��6�7�8�9�>���x@�2 @.� TRQ��$%f��4ր����_U����z��Oc <� �����Ȩ3�2��LL�ECM�-�MULTIV4�"$��A
2q�CHILD>�
1���z@T_1b  4� STY2�b4�=@�)24����@��� |9$��T��A�I`�E��eTOt���E��EXT����ᗑ�B��22(�0>��@��1b�.'��}!�A�K�  �"K�/%�a��R���N?s��=�O�!M���;A�֗�M�� 	��  =�I�" �L�0[�� R�pA��$JOBB�����ނ�TRIGI�# dӀ����R�-'r0��A�ҧ��_M��b7$ tӀFL6�BsNG�A��TBA�  ϑ�!��
/1�À�0���R0�P/p ����%�|��Bqh@W�
2JW�_RH��CZJZ�_zJ
?�D/5C�	�ӧ�t�@��Rd&�������ȯ�qGӨg@N�HANC��$LG /��a2qӐ� ـ@��!A�p� ���aR��0>$x��?#DB�?#3RA�c?#AZt@�(p.�����`FCT��ƕ�_F࠳`�SM��!I�+lA�%` � ` ���$/�/����[�a��M�0\��`l��أHK��AEs@�͐�!�"W��N� SbXYZW�`�"�����6��C����'/  . II��2��(p�STD_Cp�t�1Q��USTڒ�U�)#�0U[�%�?IO1��� _8Up�q�* \��=�#AORzs8Bp;�]���`O6  RSY�G �0�q^EUp��H`G�� ���]�DBPXWO�RK�+* $S�KP_�p�ÍA�T}R�p , �=@�`����Z m�OD3��a _C"�;b�C� �GPL:c�a�tőS�D�W�3Bb�����P��P )D�B�!�-�B APR¼�
I�Ja3��. �/�u����� �LBuY/�_�S��0�_^���PC�1�_�����~�EG�]� c2�_�SVPRE.���R3H $Cއ�.$L8c/$puSނz IkINE�fWA_D1%�ROyp �������q�c7 t@�fPA���RET�URN�b�MMR�"U��I�CRg`E�WM@�SIGN�Z�A ���e� �0$P'�1$�P� ��2p�p't��+pD�@ �'��bdNa)r�GO_A�W ��@ؑB1fI�CSd�(�CYI�	4���`1w�qu��t2�z2�vN�}���E}sDEVIs` 5 P $��SRB��I�wPk��I_BY���"�yT7Q�tHNDG�Q6 H4��1�w�>�$DSBLC�ào��vg@��|tL��a7O�f@]���FB���FEra8�ׂ�t}s���8> i�T1?���MCS���fD �ւ[2H� W��EE����%F����t����9� T�p��x�NK_QN:�����U��L�wKHA�vZ' ~�2����P~r�q7: �N=MDLn���9�� ��ٱh����!e����J��~�+���� ,�N�D����3��Ւ8G!aqSLAd�7w;  ��INP���"�����}q_ �4<j�06`C� NU��W  D�Lק��SSH!�7=M��q���ܢӢ����g���>P +$ ٰ�٢��^��^�Y�FI B\��Ă���'A	'AWl�N�TV��]�V~�X�SKI�#T���a�ۺ$�T1J�3:3_�P��SAFN���_S}V�EXCLU��*N@�DV@Ll @��Y����S�HI_V�
0\2PPLYPR�o�HIM�T�n�_M�LX��pVRFY�_�Cl�M��IOC�UC_� ����O�q�LS�0v�FT%4Q�����@�P�E$�t��A��CNFt�6եu��p��4ACHD�o����6��AFC CPlV��TQTP?�� �� ?`�@TA�@�0L@� ��N��]� �@����T��T! �S����te@{RA qDO�� w2��&�!n��_1�#�H!�̔�΀K��B|�2��MARGI��$����A ��_�SGNE�C;
$ �`�aqR0��3��@� B��B��ANNUN�P?���uCN@�`%0����� ���BEFc@I�RD� @Q�F���4OT�`�sFT�HR,Q�ŴCQ0�M��NI|RE������AW���D{AY=CLOAD�t�;T|�<S5}�EFF�_AXI��F`d1QO3O��Eq��@__RTRQE�G�Y���0RQj�!Evp ���F�0f��R0 �t �AM�P�E<� H 0�`œ^�`Ds��DU�`���BCANr� I?�`N �ErIDLE_PW�RI\V!n0V�wV�_[ ꐅ �DIA�G�5J� 1$-V�`SE�3TQl��e��Pl�^E�_��j�VE� �0SWH�q(� �bd�Gn�OHfxPPHk�IRAl�B�@�[��a�bk� �w3�O � ��v���I�0 �pR7QDW�MS-�%�AX{6j�LIFAE�@�&�MQy�NH! Q%��F#C����QCB0�mpN$�Y @ΟaFLAl���OV�0]&HE��l�SU'PPO�@u�y��@1_�$��!_X83�$gq�'Z�*W�*B1�'0T�#`�k2XZáj�+Y2D8CY`T@�`BN����f� ��C�k���ICTA��K `�pCACH��ӫ�3����I��bN�ӰUFFI� @\��@��;T��<S6CQ�.�MSW�5L 8�	�KEYIMAG�cTMLa��*Ax�&E����B��OCVIE�R-aM ��BG�L����y�?� 	���П4N�:�ST�!�BP�D,P��D��D��@EMA�I䐔a��s�FAUL|RObB�c�� "spUʰMA"`T'`E�?P< $S��S[ � ITw�BU!F�7y��7�tN[�L'SUB1T�Cx�o�8R�tRSAV|U>R�'c2�\�WT���P �T�*`Sn�_1PbU����YOT�bK��P«�M��d���WAX���2��X1P��S_uGH#
��YN_�.��Q <Q�D��0����M�� T��F�`|�\�DI��EDT_Pɰ:�IR��b�GRQM�&��HJq�a���׀��Fs�� S (�SV qpB��4�_�.��a��?T� �@����B�SC_R]1IK >B'r��$t��R"A#u��H�aDSP:FrP�lyIM|Sas�qzՄ�a� U>w� <1%sM�@IP��s��0`tCTHb0ЃTr��T`�asHS�cCsBSCʴq0� V�����S��_D��CONV�E�G���b0^v1PF�Hy�dCs�`&a?ASqC���sMERg�>�aFBCMPg��`�ET[� UBFMU� DU%P�D�:12�CDWy�p�P�C�G�[@NO6�:�V � ��� ���P���EC�����w��A���`��WH *�LƠ�Cc�W���� Y�賂��р�q�|񠀖��A��7}�8B}�9}�H ���1��U1��1��1��1ʚU1ך1�1�2���2����2��2��2���2ʚ2ך2�2*�3��3��3����U3��3��3ʚ3ך�3�3�4��QEXT[�X[b�H``@t&``z�k`˷$����FDR�YTPV��RK"	��K"�REM*F��]"O�VM:s/�A8�TR�OV8�DT�PX�MXg�IN8ɉ W��'INDv�["
�ȕ`K ^`G1a�a��@Q%r7Da�RIV���u"]"GEAR:qI%O.K(�[$N�`����,(�F@� \#Z_�MCM<0K! �Fr� UT���Z ,��TQ? b�y@\t�G?t�E �|�.�>Q����[ j�Pa� RI�E���UP2_ 3\ �@=STD	p<TT���������a>RwBACUb] T��>R�d)�j%C�E��0��IFI��0��i��{�4�PTT��FL{UI�D^ �?0gHPUR�gQ�"�r��a�4P+ I�$���Sd�?x��J�`CO�P�SVRT|��N�x$SHO* ��CASS��Qw%�pٴBG_%��3�����FO�RC�B��o�DAT�A��_�BFU_�1��bb�2�en�b0��`� |��NAV	`S������$�S�B~u#$VISI��6�2SC	dSE����j�V��O�$&��BK�� ��$P�O��I��F�MR2��a ��	��`#ǀ�&�8�O� (�_r����+IT_^��ۄ)M�����DG�CLF�DGDY&�LD����5Y&�ϤQ$Y�M됇CbN@~{	 T�FS�P�Dc P��W�cK $EX_WnW�1%`]��"X3�5��G+�d ����SWeUO�D�EBUG��-�G�R��;@U�BKUv��O1R� _ PO_ )������M��LOOc>!S�M� E�R�a��u _?E e >@�G�TERM`%f>i'�ORI�ae 9gi&�`SM_�`>RBe hi%V�(ii%�3UP\Bj� -���e��w#� �f��G�*ELT�O�A�bF�FIG��2�a_���@�$�$g�$UFR�b$`�1R0օ� OT_7�F�TA�p q3NST�`PAT�q�0�2OPTHJ�ԀE�@:�c3ART�P'5p�Q�B�aREL�:�aSHFT�r�a�1��8_��R��у�& � $�'@i�
�����s@bSHI�0�Uzy� �QAYLO�p �Oaq�����1����pERV��XA��H ��m7�`�2%�P�E3��P�RC���ASY1M�a��aWJ07�����E�ӷ1�I��ׁU�T�`Oa�5�F�5P��su@J�7FOR�`ML P�GRO!k]���5&�0L0���HOL ;l �s2T����OC1!E�$OP��qn���#$�����$��P�R^��aOU��3e��R�5e�X�1 ��e$PWR��IMe�BR_�S�4�� �3�aUD���`�Q�d]m��$H�e!�`�ADDR˶HR!G �2�a�a�aQ�R��[�n H��S����%���e3��e���e��SE���L�HS�MNu�o���Pªq��0OL�s߰`ڵ<�I ACRO��&1��ND_C�s��A<fdK�ROUP��R!_�В� �Q1|�= �s���y%��y-��x�� �y���y>�=A�����AVED�w-��ux�`(qp $_���P_D�� ��'rP�RM_��HT�TP_�H[�q (ÀOBJ��b �$˶LE~3�P��>\�r � ����J��_��TE#ԂS�P�IC��KRLPiHI�TCOU�!��L ���PԂ������PR���PSSB�{�JQUERY_FLAvs��@_WEBSOC����HW�#1��s��`<PINCPU(���O���g������d��t��O��IwOLN�t 8��yR��$SL!�$INPUT_&U!$`��Pw�֐SL.���u����2�.��C��B�I�Oa�F_AS=v�$L+ਇ+�A��bb41�����Z@HYʷ����#qe�wUOP:w `v� ϡ˶�¡�������"`PIC`���� �	�>H�IP_ME��v�7x Xv�IP�`(��R�_N�p�d��`�Rʳp�ױQrSP �z�C��BG(� ��9M�Av�y lv@C�TApB��AL TI��3UfP_ ۵�0PS6ڶBU_ ID� 
�pL � `�pr��L��0z)�����ϴ�NN�_ O��I�RCA_CNf� �{ �Ɖ-�CYpEA������� �IC�ǫ�tpR�=Q�DAY_
��NTVA�����!��5�����SCAj@��CL��
����
���v�|`5�VĬ2b�l�N_�PACV�n�
���w�})� T��S�����
��e����T� 2| ��� �v�~��֣�ذLAB1��_ �חUNIX��ӑ I�TY裪��e���p�� ��<)���R�_URL���$A;qEN ���s`vs�TeqT_U���iJ��X�M�$���E�ᒐR祪�� A��,���JH���FL�y��= 
���
�wUJR|U� ���AF�6G��K7��D>��$J7�s��J8B*�7���3�E�7���&�8\�)�APHI�Q4�y�DkJ�7J8R��L_K�E'�  �K�͐LMX� � �<U�XRi�����WATCH_VAZqxu@AំFIEL`�b�cyn���:� � bu1VbwPCTX�j�;�LGE�߄� !��LG_SIZ΄�[8XZm�ZFDeIY p1!gXb ZW �S `�8�m��� ��b ��A�0_i0_�CMc3#�*'F Q1KW d(V(Bbpo pm�p� |Io�1 p�b pW RS��0 7 (C�LN�R��۠�DE6E�3����c�i���PL�#�DAU"%EA`q�͐�T8". GH�R���y�BOO�a��� C��F�IT0V�l$A0��RE���(GSCRX����D&�|ǒ�qMARGI4� Sp�,����T�"�y�	S��x�W�$y�$���JGM7MNCHLt�y�FN��6K@7�r�>9UFL87@L8F�WDL8HL�9STPL:VL8"�L8s L8�RS�9HOPh;��C�9D�3R��}P�'IU h�`4�'�5$ ��S2G09�pPOWG�:�%`�3,64��N9EX��TUI>5I� �ӌ������C3�C<0'�@,�o:��&�@�!Naq�vcANAy��Q�A�I]�gt7Ӝ�DCS����cRS�cRROXXO"dWS�ÂRoXS{X�(IGNp 
Ђ=10 ܰ�[TDEV�7LLB��; B��C �	 8�Tr$f/蛒h����3A�a�	 �W�萦�Oqs�S1Je2Je3Ja��BSPC � �ƋG`-T��%��Q�T�r@X�&E�fST�R9 �YBr�a �$E�fC�k�g��f	v89�CB� L���� � ��u�xs뀔�g�q��jt��!�#_ ����ʐv�#Ӡ �s ��MC�� ����CLDP᠜�TRQLI ���y�t�FL���rQ��s5�D���w~�LD�u�t�u�ORG���1�RESERV��M����M�Œ�t��� �� 	�u�5�t�uSVH��p��	1�����RCLMC��M�_��ωА��_C�MD�BGh�I����$�DEBUGMASP������U�$T8P���EF�d��pFR�QҤ� � ~K	HRS_RU4��bq��A��$EFR3EQ6u!$0YOVER�k��f��PU1EFI�!%Gq�� �7�
Y�z�ǐ \����E�$9U�`��?��
�SPSI`��	��CA ���ʲ�σUY�%��?( 	��MIS�C�� d��aR5Q��	��TB� �c ���A��AX����𑧪�EXCESHg�9d�M�H�9�au���}qd�SC�`� � H�х�_������������pK�E��+�� &�B_^, FLICBtB� �QUIRE CMO�t�O��얩qLdpMD� �p{!��5�b���$L�MND!��I����L� �D;
$INAU9T�!
$RSM���PN�b�C����PSTLH� 4nU�LOC�fRI"�v�eEX��ANG.R�.���ODA]��bq��� �RMF0 ����icr�@mu����$�SUPiu��FX��IGG! � ���cs��#cs
F ct��ޒ�b5��`E��`�T�5�tC��g�TI���7�M���� Mt�MD���)��XP��ԁ��H��.���GDIAa��Ӻ�W�!P��0af���D@#)�Ҹ�㥀��� �C�Up V	���.���Or�!_��� �{`0�c������ |�P|��0� ��P{�KqEB��e-$B��o�=pND2ւ�����2_TXltXTR�AXS������LO�: ����}�L����C�.�&�[�R�R2h��� -��!A�� d$OCALI���GFQ:j�2F`RINbn�w<$Rx�SW0ۄܨ��ABC��D_�J��{�q��_J3:��
��1SP, �q�P����3��H�9p
q�#J�3n����O�QIM耯�CS�KP�zb7?SbJ+ᯂQb�y�����_AZ��/�E�L�Q.ցOCMP0�ð�� RTE��� �1�0 ���1���@ ZSMG��0�Э�JG�pSCyLʠ��SPH_�P���f��q�u�R'TER��n�Pk�)_EP�q�`A� �c̯��DI�Q23=UdDF  ����LW�VEL�qIqNxr�@�_BLXP.��Y/�J��'>$  �IN���B]�C�9%�".�8!:6p_T� �F%a"�"p^$��k)�~p�DHʠ��\�9`�$Vw��_�A$�=��~�&A$���S�h��H ��$BEL� m��_oACCE� 	8<�0IRC_�q��@�NT��c$SPSʠ�rL��� M4�s9 .7��GP/6��9�7$3�73S2T�͡_Ga�"�0�1��8�17_MG}�DD�1�~�FW�p��3�5$3�2�8DEKPPA�BN[7ROgEE �2KaBO�p�Ka���1�$USE_tv�SP��CTRT�Y4@� �� <qYN�g�A�@�FR �ѢAM:�N�=R�0O�v1�DINC(��B�4����GY��ENC�L���.�K12��H0IN¿bIS28U��ONT|�%NT23_�~�fSLO�~�|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1����PERCH  �S��� �W���SlщR ��l����E�0�0P	AS2EeL�DP7�O�NUЉZ�f�VTRK�RqAY"�?c��a S2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gBT��DUX �2S_BC?KLSH_CS2Fu :��V���C-�esRoz|�A�CLALMJTp@��`� �uCHKe |����GLRTYp� ��8T��5���_�ùT'_UM3��vC3��1�Z���LMT��_ALG��%���0�E*� K�=�)�@5F�@8 9��Nb��)hPC�Q)hHpТ��5�uCMC��\�0�7CN_��N��L�;SF�!iV�B���.W���S2/�ĈCAT�~SH�Å��4  V�q/q/V�T1�f�0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e��R� @B�_Wu�d@�!a��#`��#`�Ih�Iv�I�#F��S�:X��I�0VC00��֢1ܮ�0�⦇JRKܬ!��<�D�BXMt�<�M�_sDL�!_bGRVg�``��#`��#A�H_%�8?��0��COS��� ��LN#���ߥŴ�  ��=������꼰�<�1Z���VA�MYǱ:���᯻[�THET=0�UNK23�#��l�#ȰCB��CB�#Cz�AS�ѯ����#����SB�#��'GTSkZAC�����&���$DU�phg6�j��E�%eQ%a_��x�NEhs1K�t�� y��A}Ŧկ׍�����LCPH����^U��Sߥ ����������!��(Ʀ�V��V�غ ��UV��V��V
�V�UV&�V4�VB�H��@������d�����H
�UH�H&�H4�HB�O��O��Os���O���O��O
�O�O*&�O4�O(�F�Ҫ��	���SPBA?LANCE_J�6�LE��H_}�SP�>!۶^�^��PFULCb�q����K*1�UTO_<�p�uT1T2�	
22N�q2VP�M�a�� i�Z23	qTu`O��1Q�INSEG2�QREV�PGQgDIF�ep)1�U6�1��`OBK�q�j�w2,�VP�qI�L�CHWAR4B�BA�B��u$MEC�H��J��A��vAX��aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ�@��C1_ɒT �� x $WEgIGH�@�`$��d\#��I�A�PIFvAN�0LAG�B��S�B�:�BBIL�%OD��`�Ps"ST0s"P:�pt � N�C!L ��P 
P2�Aɑ � 2��Tx&DEB�U�#L|0�"5�M'MY9C59N��$4Ώ`$D|1 a$�0ېl� > D�O_:0AK!� <@_ �&� �q�A��B�"�� NJS�8_�P�@���"O�p ��� %�T7P?Q�TxL4F0TICK�#�T1N0%�3=p�0!N�P� u3�PR\p�A��5��5U0PRO�MP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a�@�RU�COD�#FU�@�&ID_�P�E8�2B> G_SUFF��� �#�AXA�2DO�7/�5� �6GR�#��DC�D���E��E-��DU4� ��_ H_FI�!�9GSORD�! R 236s�HR�AN0�$ZDT�El.�p�!X5�4 *WL_NA�1�0�R>�5DEF_I�X�R F�T�5�"�6�$�6�S�5�UFISm�#�m1|��40c�3�T6�44􁆂�"D� ?rfd��#D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D �S�D�U�D>b�B�c�E �S�Dd�B�&2v2a�C �ʑ�E�R�E�S�C9wwu�H�0P} d�0,aĂ�F0W�h�u�cR�VI�TE�qY4�� �!LOM�B_�r�w0s"VI]S��ITYs"Aۑ}O�#A_FRI���~SI,a�n�R��07��07�3�#s"WB�W�Q��%�_���AEAS{#�B��P|�x`WB8�45�55��6|#ORMULA�_I���G�W�� h 
>75C?OEFF_O�1&H)��1��Go�{#S� �52CA� :?L3�!G�Rm� � � �$�`�v2X�0TM�g���e�2�c��3�ERIT�d�T� ��  �LL�Dp`SΛ�_SVkd��$��v� �.���� � ���SETU,cMEAG@�@Πt �!HR>L � � (�  0��l��l��aDw��R�0�a�a}d�]�d��B��Ay`�Gax`��[Ѐk@R�EC[Qq�R0MS�K_A y�� P~_!1_USER������*���VE�L����-�!��I�zPB�MT�1CF}G���  �0z]O�NOREJ �0l���[�� �4 e���"�X�YZ<SB� 3�Iށ�_ERRK!� U ѐ�1�@c�Ȱ�!��>�B0BUFI�NDX��R0� MO�Ry�� H_ CU ȱ�1��dAyQ?�I�>Q$ +��a����� \�G{�� � $SI�0h��@2	�VOv�qО- OBJE| w�A�DJUF2yĈ�AYh�����D��OUKPp����AMR=��T��-���X2DI�R����Xf�1  D#YNt�0�-�T� ���R��0� ���OP�WOR�� �},B0SYSBU����SOPo���zډUy�XP�`K���P�A�q������OP
�@U���}�"1^��IMAG۱_ ��п"IM.���IN�������RGOVR!D"ё�	���P����@  >gplcC��L�`�BŰ?l�PMC_QE�P�1N��Mr��1212R�"�SL�| ��� �R OV�SL=S�rDEX�\a`��2�:�_ "���P#���P������2�C �P>���#�_ZERl�8��:���� @��:��O�PRIy��
�[�g@e���s�P�PL����  $FWREEY�EU�~�TZ��L����T��� ATUSk�,1C#_T�����B�������p�Vc1��P���C Dc1�к���LQ�����MQ��ۡL�XE@��x�5IP�W��` ��UP��H`&aP!X;@��43�����PGY��g�$SUB���q�����JMPWAIT8~ ���LOW���1wē CVF_A�0�b�R�Z��CC ��R$��28IGNR�_PL��DBTB2� P*a�BW@.2t�U�0-IG��!@=I�TNLN,��RBѡb�N!@��P�EED~ ��HADCOW� ��t���E��p����PSPD��� L_ A�нP���	#UNq � �RP (�LYwPa��}��PH_PK����b�RETRIE���x���2�R!D@FI��� ���V �$� 2�d�DBG�LV<LOGSIYZz�baKTU��r�$D��_TXV�EM�Cڡ)�� �-�R�#�r��CHECAKz����L���ϰ�q)�L��NP�A�`TJ"����)1P4����
�AR�"�BC =Sa��O�@����ATTS�u䡳&� 0w�^a�3-#UX^�4��PL�@Z�� $�d��qSWITCH��h�W��AS���f�3LLB���� $BA�Dvc��BAMi��6I��(@J5��N�UB�6[F
A_KNOWhK3qB"�U��AD+H�c� D��IPAYGLOAq�9p�C_����GrѼGZ�CLqA�j��PLCL_6� !4��BOA?�T*7�VFYCӐ�J(p��D�I�HRՐ�G$�TB��6�J(�zQ�_J�A �B�AN�D����T�BQ������PL@AL_ ��0 =�TATe��pC��D�CE����J3�P�V� T�PDCK^�)b���COM�_ALPH�ScBE<�߁�_�\��X�x\� �s ���OD_1�J52�DDM�AR<�h��e�f�cQ�TIA4�i5�i6��MOM�(��c�c�c�c�cV�B� AD�cv�cv�cPUBP�R�d<u�c�<u�b}"�1���� L$PI$��pc@��G�y��I�yI�{I�{I�s�`�A���v��v�J�b��a��HIG�3�� �0���5�0�f��?�5N�5�SAMPD Ƣ�0����;@�S ��с6��� 1���� ���`���`�1�K�P��`腽P�H��IN1��P��8� T�/��:�z�Q�z���/GAMM&�S��$GET������D^d>�
$�PIB�R��I��$HIB��_���1��E=�b�A�9�*�LW� W�N�9�{�*�Zb��:�QCdCHK0�j�ݠnI_��M�J� �Roh�Q ��sJ�-v|��S �$�X� 1�N�I�R�CH_D$R1N���^�LE���i�p�Zh8�ţMS�WFL/M�PSC�R�75�Ҽ ��3 �"Ķ�6��`��ع��紙��0SV���P'������GRO<�g�S_SA=AH�,=ńNO^`Ci� _d=��no�O�O�x������p�B�u�ȐcDO�A��!�ں�*� t�:�Z1f�;�7����C�FMmu� � F�YL�snQ ��@� ���"��<s�	�Ҁ���nQ૰<3M_Wl�����\p��(�o�MC��P���Q�����hpM.�pr� ��!��$��WM��ANGL �!�AM�6dK�=dK�DdK��TT7�Nk@��3��#�PXC OEc�QZp��hp	nt� ���OM���ϑϣ� �����`� c�Z0es^a_�2� |a�J� �i���c���cJ��j��0���jA� �Qy�>��  �@{��P�1�PMON_�QU�� � 8�60QCOU��Q�THxHO��B H�YS�0ESPBB U�E- 3�f0O�4� � c P�^�RU�N_TO��I�O��� P�@���INDE�#_PG�RA���0��2��N�E_NO��ITxf��o INFO���a"�����H�O�I� (*�SLEQ!�*�*�Q �OS��l4� 4�60ENABy� PTION�3��r���^GCF�!� �@60J�Q���R�d!��erP�EDIT�� ��� ��KAQ"� �E�(�NU'(AUT<Y�%COPYAQ�(2,�qe�M�N< @+^��PRUTm� C"�N�OU�2$G���$RGADJZ��u2X_��IX�P���&���&W�(P�(�~��&9�� 
�N�P_�CYCy�e1RG�NSc�{�s�LG�O£�NYQ_FREQSrW@��X1�4�L�@�2P0�!�c@�"�CRE��Mà�IF�q�NA���%�4_Gf�STA�TU~�f��MAI�L��|CIq�=LA�ST�1a*4ELE�Mg� ��QrFEASIt;�ւΰ ��B"�F�AF����I� ��O2�E u�&vBAB��PE� =��VA�FzQ�I��TqU�[��R��S�FRMS_TRpC�Qc���C��Z�
��1�D XI�,2ns؆�	MB? 2� `��� N�3V�R2WR*����p�R^W�wj�DOU�2^�N�,2PR`�h=�1GRID��oBARS!�TYu�Z�Op�� �|_�4!� �R�TO|��d� � ����POR�c~vb�SRV�0)"dfDI[�T�`;aNd�pXgD
�Xg4Vi��Xg6Vi%7Vi8:av�Fʒg��z $VALU��C0�3D1AC�ad�� !pf���S1�1-ȆAN/��c��0R�]11ATOTcAL����=sPWE3�I�QStREGENQzfr��X�H�]5	�v( TR�CS�Qq_!S3��wfp�V�!��r��BE�3�PG0B��( sV_H�PDqA(��p�S_Ya����i6S��AR(�2�� �"IG_S!E�3�pb�5_� �t{C_�V$CMPl��DEp�G���IBšZ~�X�
��Fm��HANC.� �p Qr�2���I#NT9`cq�F����MASK�3�@OVRMP �PD�1-� �W�QaХT�l�_�RF�{�V�PSLGP�g�9�j5���,�;pDpS���4��cU��.�}�TE����`���`k���Jx^�Y�y3IL_Mx40�s��p��TQ( �P��@����V.�C<��P_ �R�F�M]�V�1\�V1j�2y�2�j�3y�3j�4y�4 j���p۲������vܲIN�VIB8�P6�#��*�2&�22�U3&�32�4&�42���6���SJ�  ��T $MC_F,K `� �L>�J�х1pMj�Iу��zS� ��1���KE�EP_HNADD"��!鴓@�C��0A	��Q����
�O!��v ���p
�և
�REM!�	�Cq�RF��]�b�U�4e	�HP�WD  �S�BM���PCOLL�AB*�p��/q�2�IT/0��Q"NO1�FCALp⎵��7� , �FLv�A�$SYN���M���Ck��RpUP_�DLY��zDE�LA9�Dq�2Y A�D(�3��QSK;IPO�� �`� �O��NT����c�P_� ��׾ ��cp�� �q�ٞ��o`��|`�� �`�ږ`�ڣ`�ڰ`��=9�!�J2R0  �lX�@TR3H�� 1AH� �H���$ �RDCq��� �� R�R, 5��R��1��E��5TRGEp�_C��RFLG"����W�5TSPC��1UM_H��2/TH2N}Q�;�� 1� ��;��Q02 � D� ˈ��@2_PC�3W�S���1Y0L10_Cw2x�-���7 � $\�  U@��V7�����0��VU\����� rd��C *��7��DZ Gs�RUV�L1[�1h���10]�_DS�������PK 11�� l�ڰ����q��AT ?��$�Q[7�� ���K 5T���HOMME� ��c2h�n�����&0
`3h���!L3E *�c4h�hz�����5h���	//-/�?/ �`6h��b/t/�/�/�/�/�7h��/�/??'?9?
�8h�\?n?�?�?,�?�? _S����  �Aa{p���_�]�Ed� aT=�nD4vnCIO�ҎII@`�O��_O�P�E�C.rfBXPO{WE	�� X@��f��$$�Cd�S�����4�A3�3� �@�sSI��GP�0�QIRTU�AL�O
QAAVM_WRK 2 7U� ?0  �5Qn_rzXk_�] �\A	�P�]�_3�8P��_�_�Ve�\#m/o�Q`5ojo|o�dHPBS��� 1Y� <Xo�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯz�bC$�AXLM�@tiAQ��c  d��IN����PRE�
�E�J�-�_U�P��[�7QHPIO�CNV_�� �	�Pr�US>��g�c{IO)�V 1U[P $E`��Qս9lҿ8P?��i@��� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o��o�m�LARMRECOV a���-���LMDG ���ɰ�LM?_IF ��� ை����zv����%�6�, 
 6�_��r漅�������̍$w���׏���8�J�\�n����NGTOL  a�� 	 A   ���ț�PPINFoO ={ <v�����1��   I�3�a�"rP���t��� �����ί���>�o����j�|������� Ŀֿ�����0�B��PzPPLICAT�ION ?����J��Handling�Tool �� �
V9.30P/�04ǐM�
88g340�å�F0����202�ťʚϬ�7DF3��M̎��NoneM�F{RAM� 6���Z�_ACTIVE��b  sï�  ~p�UTOMODz��A���m�CHGAoPONL�� ���OUPLED 1ey� �������g�CUREQ �1	e{  T�
��	p��w����#r���e�HN���{�HTTHKY��
$r��\[�m���� O�	�'�-�?�Q�c�u� ������������ #);M_q�� ����% 7I[m��� /���/!/3/E/ W/i/{/�/�/�/?�/ �/�/??/?A?S?e? w?�?�?�?O�?�?�? OO+O=OOOaOsO�O �O�O_�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_oo#o5o GoYoko}o�o�o�o�o �o�o1CU gy������ �	��-�?�Q�c���1�TO��|�p�DO_CLEAN��|n��NM  �� �B�T�f�x����%�DSPDRY�R��m�HI���@ /�����,�>�P�b��t���������ίj�MAXa�ۄ��������Xۄ������p�PL�UGG��܇�ӌ�P�RC��B� ���ׯF�OK���ȔSEGF��K������ �.�����,�>�v���LAPӟ澨�� �϶����������"��4�F�X�j߯�TOT�AL�7���USE+NUӰ�� �������1�RGDISPWMMC����C��&��@@Ȓ��Oѐ������_STRI�NG 1
��
��M��Sl��
A�_ITEM1K�  nl�g�y�� �����������	�� -�?�Q�c�u����������I/O S�IGNALE��Tryout M�odeL�Inp���Simulat{edP�OutOVERRА� = 100O�In cycl�P�Prog A�borP���S�tatusN�	H�eartbeat�J�MH Fauyl��Aler�	 ������*8<N` ׃G� ׁY�c����� ////A/S/e/w/�/��/�/�/�/�/�/wWOR��G�-1�?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO8�O�O�NPOE� �@E;�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo�BDEV�Nu`�Obo�o �o�o�o�o�o, >Pbt��������PALT ��E?�A�S�e�w� ��������я���� �+�=�O�a�s����GRI�G뽑1��� ���	��-�?�Q�c� u���������ϯ�� ��)�����R�a� ՟;���������ѿ� ����+�=�O�a�s���ϗϩϻ���O�PREG��y���-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_��q����$ARG_�-0D ?	������� � 	$��	+[��]����������SBN_CONGFIG���� ��CII_S?AVE  ��)����TCELLSETUP ���%  OME_I�O����%MOV�_Hn�����REP�d�����UTOBA�CKY���#��FRA:\�� �����)�'`l ���&� 7"�� 24/0�6{  09:35:24�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� ,,		�����O�G�O __#_%_7_q_[_�_ _�_�_�_�_�_�_%o����D�@TSK � �M&,O��UP3DT�@EGd�`�F�XWZD_ENB8ED��fSTADE��ܖe��XIS�UNOT 2��&�(��� 	 0|�} Z�0&�? �<_ �/� K��pp�T<�bp�p�8t�}V��)q{|��t�� B=|�o���;9Յ�!{D�x�Q\��gMETc�2Lf�E� P qA|h�iA��A��B-��B��B�y��}?y�J�?��?:��&@5�W?U��s@���}S�CRDCFG 1��� ��z�����ԏ�����Q=���H�Z� l�~�����	�Ɵ-�� ��� �2�D���域���GR�`�`�O���0kNA����	��n��_EDC@1n��� 
 �%-�0EDT-q����L%�p��"���-������������^��  ����2����*�R�bB���*� q���ϧ���3bϮ� @Ͻϯd?�����=�O���sϏ�4.ߞ�{��� ��W���	�߱�?ߏ�5��j�G����#�� ����}�6��6� �Z�����Z����I��7�����&��΀��&m������8^ҿ����	͇� 9K�o��9*�w��	�S��;��CR����B/ T//�/��w//���РNO_DEL�����GE_UNU�SE���IGAL�LOW 1���2p(*SYS�TEM*�s	$SERV_GR�;�B0�@REGK5$8m3�|B0NUMp:�3��=PMU� �u�LAY�p�|?PMPALD@�5�CYC10�.�>x�0�>CULSU�?0�=�2�AM3LOWD�BOXORIt5C�UR_D@�=PM�CNV�6D@1�0�>�@T4DLI��`=O_9	*PRO�GRAJ4PG�_MI�>�OPAL(�E_UPB7_B>�$FLUI_RESU�7p_z?�_�T#MRY>h0�,�/�b �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� ��������"�LAL_OUT �1;l���WD_�ABOR�0?d�I�TR_RTN  �����g�NONgSTOǠ�� 8�CE_RIA_IL0��ۀ��ŀFCFG ��x۔��_LIMY2�2ګ �  �� 	i�J��<�e�g��5��  9��������
����u��PAQPGP ;1�����Q�c�u�4�CK0����+C1��9��@���P�C��CV��]��d
��l��s��P����C[٤m��v���������� C�j���-���?�Â{HE� ONFI�P�q�G�G_P�@1� �%��������ǿٿ����G�KoPAUSaA1�ۃ �B�W��E� ��iϓϹϟ������� ���#�I�/�m��e�����M��NFO �1"��� �7��ߖ��C w��Bb?	�;���8����,,�MA�@�� �ģ�C�Tp���1VC3�����"��3��h3�E�ŀO����c�COLLECT_�"�[�����EN�@��y���k�N[DE��"�3��"1234567890��\1��H ��֕H&��)M� r�\,L�^���]+���� ��������C 2 �Vhz���� ��
c.@R �v���������� ����I�O !���q����u/�/�/�/C'TR��2"'-(׀^)
��.R�#R-�*W�^ 9_MOR�$� �;�l5��l9�?r?��?�?�?�;E2��%JS=,W�?@�@��CR׀K)DցC�R��&u�XOWAWBC4 � A&��׀x׀}A"@Cz  B�@�CG�B8��AC � %��׀ց:�d�43 <#�
�E���I�O�C=A�I��'GM?�C�(�S=���Qd=AT_D�EFPROG ��;%�/m_APIN�USE�V�ۅ�TK�EY_TBL  �s�ہ���	
��� !"#$�%&'()*+,�-./�:;<=�>?@ABCDPG�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������Ga��͓���������������������������������耇����������������������!�PLC�K�\���P�PSTA�n��T_AUTO_�DO��NFsIN�D���n��R_T1wT2N����5�ŀTRLCPLET�E���z_SCR�EEN �_kcscÂU���MMENU 1)O� <�[_#�q� �,�a���>�d���t� ��ӏ����	����� Q�(�:���^�p����� ��̟�ܟ�;��$� q�H�Z���������� Ưد%����4�m�D� V���z���ٿ��¿� !���
�W�.�@ύ�d� vϜ��ϬϾ������ A��*�P߉�`�r߿� �ߨ��������=�� &�s�J�\������������'�,�p_M�ANUAL�EqD�B
12�v�iDBG�_ERRLIP*�{h! 0��������g�NUMLI�M�s:QOE�@DB�PXWORK 1+�{��>Pbt|��-DBTB_�qG ,��kC3!VD�!DB_AWA�Yo�h!GCP �OB=��A�_AL���o�k�Y�p�uO@�`�_�� 1-�+@
-k-6[���_M+pIS�`�@|"@�ONTIM�w��OD��&
��U;MOTNEN�D�_:RECOR�D 13�{ �<�[CG�O�f!T/ [K��/�/�/�/_(�/ �/f/?�/??Q?c?�/ ?�??�?,?�?�?O O�?;O�?_O�?�O�O �O�O(O�OLO_pO%_ 7_I_[_�O_�O�__ �_�_�_�_l_!o�_,o �_io{o�o�oo�o2o �oVo/A�oe P^�
���R ���=��a�s��� �����*�ߏN��� '���ԏ]�̏������ ��ɟ۟v���n�#����G�Y�k�}���TO�LERENC�B��0� L��g�C�SS_CNSTC�Y 24	�t���.������0� >�P�b�x��������� ο����(�:�ä�DEVICE 25ӫ ��ϟ� ������������/��AߟģHNDGDg 6ӫ� CzT�|.!ơLS 27t�S������������/�U�ŢPARAM 8Gb�A��~��RBT 2:�8�<���{CkA� ·�?  � A��8�.SB���A�?B�  ���a������.��  ����A�A�C�����c�u����C�A�D��k�p�z�A�A��HA�c ��A�	�?(uL�^p���A�Bt�/�D��C��_� 	 A=���ABffA#3�3AҊ���AY�A�Cf��a���A�J��7B]���B��Bf�fBᴠ�33Ca$.@R� (�� ���A����
/ ��//)/;/�/_/ q/�/�/�/�/�/�/�/ <??%?r?I?[?m?? �?�?�?�?�?&O8O� PObOMO�OqO�O�O�O �O�O_�OOL_#_ 5_�_Y_k_�_�_�_�_  o�_�_6oooloCo Uogo�o�o�o�o�o�o  �o	h�O�w �����
��.� 	__I'�1_�q��� �����ˏݏ��� %�r�I�[�������� ��ǟٟ&����\�3� E�W����ȯ���ׯ �"��F�1�j�E�s� ����m�������ѿ� 0���f�=�O�a�s� �ϗ��ϻ������� �'�9�Kߘ�o߁��� ��[����(��L�7� p��m������� ����$�����l�C� U���y�����������  ��	V-?�c u����
�� @+dO�s�� ������*/// `/7/I/[/m//�/�/ �/�/?�/�/?!?3? E?�?i?{?�?�?�?�? �?�?�?FO�jOUOgO �O�O�O�O�O�O__ �'O9OO=_O_�_s_ �_�_�_�_�_�_�_o Po'o9o�o]ooo�o�o �o�o�o�o:# 5��O������ ��$��H�Fz�$�DCSS_SLA�VE ;��}�w��`�?_4D  w����AR_MENU <w� >�؏���� �2�^rǏ\�n��\���SHOW 2}=w� � fr [q����Ə�����@,�>�D�b�t��� �� ��ҟϯ����)� P�M�_�q��������� ˿ݿ���:�7�I� [ς�|Ϧ��ϵ����� ����$�!�3�E�l�f� �ύߟ߱�������� ��/�V�P�z�w�� ������������ @�:�d�a�s������� ����\���*�H�N� K]o������ ��28�GY k}������ "�1/C/U/g/y/ �/��/�/�/��// ?-???Q?c?u?�/�? �?�?�/�??OO)O ;OMO_O�?�O�O�O�? �O�?�O__%_7_I_ pOm__�_�O�_�O�_ �_�_o!o3oZ_Woio {o�_�o�_�o�o�o�o Do-Se�o� �o������.�=�O���CFG >�����q��dMC:\���L%04d.CSIV\��pc�������[A ՃCH݀z�v��w�#��q����:�J�8�7���J�P�j�)�́�p�+�n�RC_OUT� ?z������a�_C_FSI� ?�� |�����@� ;�M�_���������Я ˯ݯ���%�7�`� [�m��������ǿ� ����8�3�E�Wπ� {ύϟ���������� ��/�X�S�e�wߠ� �߭߿��������0� +�=�O�x�s����� ���������'�P� K�]�o����������� ������(#5Gp k}�����  �HCUg� ������� / /-/?/h/c/u/�/�/ �/�/�/�/�/??@? ;?M?_?�?�?�?�?�? �?�?�?OO%O7O`O [OmOO�O�O�O�O�O �O�O_8_3_E_W_�_ {_�_�_�_�_�_�_o oo/oXoSoeowo�o �o�o�o�o�o�o0 +=Oxs��� ������'�P� K�]�o����������� ۏ���(�#�5�G�p� k�}�������şן � ����H�C�U�g��� ������دӯ��� � �-�?�h�c�u����� ����Ͽ�����@� ;�M�_ψσϕϧ��� ��������%�7�`� [�m�ߨߣߵ����� �����8�3�E�W�� {������������ ��/�X�S�e�w��� ������������0 +=Oxs��� ���'P K]o����� ���(/#/5/G/p/ k/}/�/�/�/�/�/ ?��/??H?C?U3�$�DCS_C_FS�O ?�����1 P [?U?�?�?�?�? �?O
OO.OWOROdO vO�O�O�O�O�O�O�O _/_*_<_N_w_r_�_ �_�_�_�_�_ooo &oOoJo\ono�o�o�o �o�o�o�o�o'"4 Foj|���� �����G�B�T� f���������׏ҏ� ����,�>�g�b�t� ��������Ο���� �?�:�L�^�������যϯʯܯg?C_RPI~>�?�;�d� _�
�}?.�p����ݿj>SL�@���9� b�]�oρϪϥϷ��� �������:�5�G�Y� ��}ߏߡ��������� ���1�Z�U�g�y� ������������	� 2�-�?�Q�z�u����� ��������
) RM_q���� ���*%7I rm����� /�ϛ�,�/W/�/ {/�/�/�/�/�/�/? ??/?X?S?e?w?�? �?�?�?�?�?�?O0O +O=OOOxOsO�O�O�O �O�O�O___'_P_ K_]_o_�_�_�_�_�_ �_�_�_(o#o5oGopo ko}o�o�o�o�o�o  �oHCUg� ������� �����NOCODE� @������PRE_CH�K B��3�A �3��< ��7��������� 	 <�����?#ۏ%� 7��[�m�G�Y����� ��ٟ�ş�!���� W�i�C�����y�ïկ ˏ������A�S�-� _���c�u���ѿ���� ���=��)�sυ� _ϩϻϕ�������� '�9���E�o�I�[ߥ� �ߑ���������#��� �Y�k�E���{�� ���������C�U� �=�����w������� ��	����?Q+u �a����� �);_qg�Y ��S����%/ �/[/m/G/�/�/}/ �/�/�/�/?!?�/E? W?1?c?�?���?�? o?�?O�?�?AOSO-O wO�OcO�O�O�O�O�O _�O+_=__I_s_M_ __�_�_�_�_�_�?�_ 'o9oo]oooIo�o�o o�o�o�o�o#�o GY3E��{� ����o�C�U� �y���e��������� ��	��-�?��K�u� O�a���������͟ ��)��1�_�q��}� ������ݯ�ɯ�%� ��1�[�5�G�����}� ǿٿ�������E� W�1�{ύ�G�u����� �������/�A��-� w߉�c߭߿ߙ����� ����+�=��a�s�M� ���ϑ������� '��3�]�7�I����� ������������� GY3}�i�� ������C /y�e���� ���-/?//c/u/ O/�/�/�/�/�/�/�/ ?)?�?_?q?K?�? �?�?�?�?�?�?O%O �?IO[O5OO�OkO}O �O�O�O�O_�O3_E_ ;?-_{_�_'_�_�_�_ �_�_�_�_/oAooeo woQo�o�o�o�o�o�o �o+7aW_i_ ��C����� '��K�]�7�i���m� �ɏۏ������� G�!�3�}���i���ş ������1�C�� g�y�S�e�������� ��ѯ�-���c�u� O�������Ͽ�ןɿ �)�ÿM�_�9�kϕ� oρ����Ϸ����� �I�#�5�ߑ�kߵ� �ߡ�������3�E� ��Q�{�U�g����� �������/�	��e� w�Q������������� ��+Oa�I ������ �K]7��m �����/�5/ G/!/k/}/se/�/�/ _/�/�/�/?1??? g?y?S?�?�?�?�?�? �?�?O-OOQOcO=O oO�O�/�/�O�O{O�O _�O_M___9_�_�_ o_�_�_�_�_oo�_ 7oIo#oUooYoko�o �o�o�o�o�O�o3E i{U���� ����/�	�S�e� ?�Q�������я㏽� ���O�a����� ��q���͟������ �9�K�%�W���[�m� ��ɯ�����ٯ�5� +�=�k�}�������� �����տ�1��=� g�A�Sϝϯω����π��������Q�c�����$DCS_S_GN CS�����#M�2�6-JUN-24 09:26 E�70��39������� X�L����������������ќM��Þ��j�����{�V�ERSION ���V4.2�.10�EFLO�GIC 1DS���  	D���X�k�X�z�M��PROG_ENB  ��b��Л�ULSE  �����M�_ACCL{IM���������WRSTJN�T����w�EM�O���ѷ�L��IN�IT EZ�O���OPT_SL �?	S�1�
 	�R575�Ӆ�7U4��6��7��5A�
��1��2��l���G�>h�TO  t���t.H�V?�DEX���d����FPAT�H A��A\�4���HCP_�CLNTID ?<+�b� l������IAG_GR�P 2JS�? �a[��D�  D��� D  B� w B�@ff�چ/B�@[��W��@�q��B��N�C�-BzBp@e`���mp3m7� 7890123�456�*�[�� � Ao�mA�j1AdA�]�
AW|�A�P�AJ-A�C/A;�A�4H���@�  �A��A�A3!_Ae�@@��B4��G ��t���
��uƨApffA�j�yAeK�A�_�AY��A�S� MC�AF��A@ �O�+/=/�O$O�c K�w(@�X�?8��@��y�/�/�/�/�/8��;d�2�5?@�~ff@x1'@�q��@kC�@�d�D@]��@Vv�6?H?Z?l?~?�8s�0l��@e�@^��@W�\)@O��@H��0?<@7K�@.V�?�?�?�?
O8_S@M00G<@�A��@<1@�5��@/l�@�(Ĝ@!�0�\NO`OrO�O�Ox'g� L_K�;_�_�__g_�_ �_�_�_o�_�_�_Yo�koIo�o�o+o�oX��"� 2�17A�@J>���R
q?�33�?Y��r��^J7'Ŭ2q63p�4�F>r��L�J@�p�Zr�
�=@�@�Qi�jq��@G Ah�@���@�T= c�<��]>*�H�>V>�3��>���J<����<�p�q�x���� �?� �C��  <(�U��; 4Vr�33��@,
���A@��?R�o D��mR�x���Q��t�� ��Z�Џ��؏�,��i�?�7N�>�(��>�@Z�=����J��G�v�G�@J�B�E�����a��@�ǐ@���@��@�Q�?L ��
�ŲI�P���&���'��@�K�����Ag�q�PC�  C���Cuy�
���ʯ ?����	�@�Գ�4���X��v����*Cz�C��8�D�h�3��6C �F�ǿB��ֿ�����E�T��� =�2�������=��^>�&$�
�Iϗ�CT_C�ONFIG K�3���e�g��STBF_TTS��
����"��������{�MAU����MSW_C5F��L  K �OCVIEW	�MI�U��㯛߭� �����������0� B�T�f�x������ ��������,�>�P� b�t������������ ����(:L^p ������  �6HZl~� �����/��KRCB�N��!� �F/{/j/�/�/�/�/��/��SBL_FA?ULT O9*^�>1GPMSK��7���TDIAG �P��U����q�UD1: 6�78901234A5q2�q���%P�� �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O �a6�I'�
�?_>��TRECPJ?\:
j4\_�7_[�?�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�O��O_ _�UMP_?OPTION��>FqTRB���9;u�PME��.Y_T�EMP  Èϓ3B����p�A�pytUNI'��ŏq�6�YN_BRK �Qt�_�EDITCOR q&qh�r_2P�ENT 1R9)�  ,&CO�LOCA_bpA_�IRVIS$r5� �&DROP_�DEFE�p_3 SO 1��cJ�2Z���J�1����L�S�EMP����� �B�ARRA_�pNO� ���&MA�IN �ESTE�IRA���&�PEG�3��&PICKUP���M�P�p 
Ж�?&SEGU������� &SU�MIRԂ�������ؓF��DA_PROENSA럝���L�� A�����1_PLACE0>�H�&
T�	��n���&ؓ�����AR����ǯy�b� ���٥�������8�J��%EMGDI_STA�u~��q��uNC_INFO� 1SI��b��������Կⷮ���1TI� ��o#����0�d�o}Ϗϡϳ� ����������1�C� U�g�yߋߝ߯����� ����Hu� �2�D�R� j�R�x�������� ������,�>�P�b� t�������������Z� �#5Ga�k} ������� 1CUgy�� ������	//-/ ?/Yc/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? ��?O%O7OQ/GOmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�?Ooo /o�_[Oeowo�o�o�o �o�o�o�o+= Oas����� �_�_��'�9�So]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�K�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�C�5� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ�������� �!�;�M�W�i�{�� ������������� /�A�S�e�w������� ��������+E� Oas����� ��'9K] o����1��� �/#/=G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?��?�?	OO5/ ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�?�_ �_oo-O#oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���_�_���� 7oA�S�e�w������� ��я�����+�=� O�a�s��������� ߟ���/�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������͟׿���� '�1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߫�ſ ���������;�M� _�q��������� ����%�7�I�[�m� ������߯������� �)�3EWi{� ������ /ASew���� �����/!+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?/��?�?�? �?/#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �?�_�_�_�_Oo-o ?oQocouo�o�o�o�o �o�o�o);M _q���_��� �	o�%�7�I�[�m� �������Ǐُ��� �!�3�E�W�i�{��� ��ß՟矝��� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}� �ߩ����������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u����߫��� ��������);M _q������ �%7I[m �������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?���? �?�?�?�OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�?�?�_�_�_�_�? �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�_� ����_�	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q��y�����˟� ۟��%�7�I�[�m� �������ǯٯ�����!�3�E�W�i��� ��$ENETMO�DE 1U��  ���������»��R�ROR_PROG %��%������TABLE  ���Q�c�uσ���SEV_NUM� ��  �������_AUT�O_ENB  �̵��ݴ_NO�� �V������ W *���������	�����+���(�:ߞ��FLTR����H�IS�Ð�����_A�LM 1W�� e����̍�+;߀��������0�?�_\����  �����²u꒰TCP_V_ER !��!���@�$EXTLOGo_REQv�������SIZ����ST�K�������T�OL  ��Dz�~��A ��_BWDU�*�Z�V�ǲ?�DID� X��Z�����[�ST�EPl�~�����OP�_DO���FAC�TORY_TUN�v�d��DR_GR�P 1Y��`�d �	p�.° �*�u���RH�B ��2 ���� �e9 ���bt�o�� �����J�5nYA���A'�q@9�u���
 JpH ��ȸo��_/��(/(B�  F!A�  @�33R"��33-@UUT�n*@P  /ȷ>u�.�>*��<���ǆ-E�� Fw@ �"�5W�%��-J��NJk��I'PKHu���IP�sF!�=��-?�  ?�/�9�<9��896C'�6<,5����-�YHv ���� �"�9d����A�FE�ATURE Z��V�ƱH�andlingT�ool �5���English �Dictiona�ry�74D St΢0ard�6�5An�alog I/O��7�7gle Sh�ift Outo �Software Update%I�matic Ba�ckup�9SAgr�ound Edi�t�0�7Camer�a�0F�?CnrR�ndImXC�Lom�mon caliOb UI�C�FnqA��@Monitor��Ktr�0Reli�ab@�8DHCP��IZata Ac�quis�CYia�gnosOA�1[o�cument V�iewe�BWua�l Check ?Safety�A�6?hanced�F�:��UsnPFr�@�7xt. DIO �@sfiRT�Wend�PErr�@LQR�]�W%s�Yr�0�P E�:�FCTN Men�u�Pv S8gTP ;In'`facNe�5�GigE`nrej@p� Mask Ex�c�Pg�WHT^`Proxy SvoT��figh-Spe�PSki�D�eJP�P�mmunicN@ons�hurE`'`_��1abconnecwt 2xncr``�stru�2z>pe�eQPJQU�4KAR�EL Cmd. �L�`ua�husRu�n-Ti�PEnv�kx(`el +R@s�P@S/W�7Lic�ense�Sn\�PB�ook(Syst�em)�:MACR�Os,�b/Offse@�uH�P8@_��pMR�@�BP^Me�chStop�at�.p6R�ui�RKj�x��P�0P@)�od@w�itch��>�EQ.<���OptmЏ>�N�`filn\=�gw~�uulti-T�`�tC�9PCM fu	nHwF�o3T�R?�f�/Regi�pr�`I��rigPFV����0N?um Selb���>�P Adju�`��x�J�tatu���
�iZ�5RDM R�obot�0sco3ve�1F�ea7��P�Freq Anl�y�gRem`��Qn��7F�R�Servo��P���8SNPX �b�rNSN^`Cl�ifQɮBLibr��3鯢0 q�����oz�ptE`ssag?���4�� -C��;��/�I_mB�MILIB�k�E�P Firmt6BU�PEcAcck@�sKTPTX_C�eln���F��1�V��orqu@imu�la�A�A�u��PAa�qU�j@�Ã&�`gev.B�.@riP�޿USB po�rt �@iP�Pa�gP��R EVNT��ϗ�nexcep�t�P��t��ſX�]VEC�Ar�b�bf�V2P�Ҧ�$����SܠS9CصV�SGEk�a��UI�;Web Pl!��ާ��Խ`�T�eQfZDT Ap�pl�d�:�ƺ� �G�ridV�playP�R�WD4�R
�.�:�n�EQ+��r-10i�A/7L*��1Gr�aphic���5d�v�SDCSJ�ck��q�5larm C�ause/��ed>�8Ascii�a���LoadnP�Up�l,�Ol�0�AGu`�6N�`���yFyc@��r�����PV��Jo��m� c�R���c����m�./�����Q�2*u:eRAJ��P�ٶ4�eqinL����8NR�T��9On�0e �Hel�HJ�`oI�a?lletiz?�H�ؘ���_�tr�[ROS Eth�q��T@�e�ׅ�!�n�%�2D�tPkg&�Upg~�(2DV�-�3D Tri�-jQEAưDefl.qEBa)pdei���� �bImπF8�f��nsp.q=��464MB DRsAMZ,#FRO5/�@ell�<�Msh�f!r/�'c%3@p,LƖ,ty@s˒xG��m��.[�� ����BU���Q�B�=ma�i�P߫�]Q����@q�6wlu����^`�xRt�?eL� Sup��`����0�P�`cr���@�R���b䚮�pr1u7est�rt~QQ��ߋL!�4O��q$��K��l Buiz7�n��APLCOO2�EVl%��CGU�O'CRG�O��DR��Of
TLS_��BU/_b��K�qN_d�TA�OxVB�_�W�ܑZ���_TCB�_�V�_�W���WF+o�V�O�W._�W�ņoTEH�o�f�O��gt�oTEj�xVF�_w�_xVGoTwB�Tw~oxVH�xVIA0��v�xVLN�yU�Mz�bo�f_xVN��xVP���^xVR�&xVS��܇ʏ��Wp��v���VGF:�L�P2_h��h�V�Hh��_g�D��h�FFo�h��g�RD�� T�UT��01:�L�2<V�L�TBGG��v�orain�UI���
%HMI���pon��m�f�"�F��&KAREL�9� �TPj��<6 SWIMESTڢF0O�<5�
"a�X� j�������ͿĿֿ� ��'��0�]�T�fϓ� �Ϝ�����������#� �,�Y�P�bߏ߆ߘ� �߼���������(� U�L�^������� ��������$�Q�H� Z���~����������� �� MDV� z������ 
I@Rv� �����/// E/</N/{/r/�/�/�/ �/�/�/???A?8? J?w?n?�?�?�?�?�? �?O�?O=O4OFOsO jO|O�O�O�O�O�O_ �O_9_0_B_o_f_x_ �_�_�_�_�_�_�_o 5o,o>okoboto�o�o �o�o�o�o�o1( :g^p���� ��� �-�$�6�c� Z�l���������Ə� ���)� �2�_�V�h� ������������ %��.�[�R�d����� ����������!�� *�W�N�`��������� ���޿���&�S� J�\ωπϒϤ϶��� ������"�O�F�X� ��|ߎߠ߲������� ���K�B�T��x� ������������ �G�>�P�}�t����� ��������C :Lyp���� ��	 ?6H ul~����� /�/;/2/D/q/h/ z/�/�/�/�/�/?�/ 
?7?.?@?m?d?v?�? �?�?�?�?�?�?O3O *O<OiO`OrO�O�O�O �O�O�O�O_/_&_8_ e_\_n_�_�_�_�_�_ �_�_�_+o"o4oaoXo jo|o�o�o�o�o�o�o �o'0]Tfx �������#� �,�Y�P�b�t����� ����������(� U�L�^�p��������� �ܟ���$�Q�H� Z�l�~��������د ��� �M�D�V�h����  Hg552}���21���R78��50��J�614��ATUP�Ͷ545͸6��VwCAM��CRIǷUIFͷ28	�N�RE��52��R6�3��SCH��DO�CV]�CSU��8�69ͷ0ضEIOuC9�4��R69���ESET���J7���R68��MAS�K��PRXY!�7.��OCO��3帨����̸3�J6˸5u3��H2�LCH�ƯOPLG�0�M�HCR��S{�MC�S�0��55ضMgDSW���OP�GMPR�M�@�0̶7PCM �R0����ض��@�51�51�<�0�PRS��6�9�FRD�FR�EQ��MCN��9=3̶SNBAE�3�/SHLB��M��M����2̶HTC�T�MIL����TPAޘ�TPTX��EL���Ѐ�8������J�95,�TUT�9�5�UEV��UE�C��UFR�VCuC��O��VIP�wCSC,�CSG8ƺr�I��WEB�H�TT�R6C�N�C�GIG��IPGmS)RC�DG��H77��6ضR8�5��R66�R7���R:�R530�6%80�2�q�J��H�6<�6,�RJح�0�4�6o64\�5n�NVD��R6�ׇR84Tg����8f�90\���J93�91� 7+���,��D0oF�CLI���CMS�� �7STY��TO�q�ژ�7�NN�OR�S��J% ��j�OL�(END��L��S�f(FVR��V3D����PBV,�AP�L��APV�CC�G�CCR|�CD��CDL@CSBnt�CSK��CT��CTBL9��U0,(Ch��y0L8C��TC �ly0�'TC(7TC���CTE\��07TEXh��0��TFd8F,(�GL8GI�8H�8Ip��E@�87�CTM,(UM�8M@8N�8PHHePL8Rd8(TSd8�W�I@VGF�GP2��P2���@�H{7�VPD�HF �VPnSGVPR�&VT��\YP��VTB7VsǋIH��VI aH'V�K��VGene �����_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/??�+?=?O?a?s?�?  H55hTp�1�1[U�3R78�<{50�9J614�9�ATU�T�4545:�<6�9VCA�D�37CRI,KUI8T�5�28-JNRE�:5�2JR63�;SC�H�9DOCV�JC\U�4869�;0�:�EIO�TsE4�:R{69JESET�;vKJ7KR68�J�MASK�9PRXuYML7�:OCO\�3�<�J)P�<3|ZJ�6�<53�JH�\L{CH\ZOPLG�;�0�ZMHCR]ZS�kMCS�<0,[5=5�:MDSW}k�[;OP�[MPR�Z�@��\0�:PCMLJR�0�k)P�:)`�[51�K51|0JPR�S[69|ZFRD�<JFREQ�:MC�N�:93�:SNByA}K�[SHLB�z�M�{�@ll2�:HT=C�:TMIL�<�J�TPA�JTPTXF�EL�z)`�K8�;��0�JJ95\JTU�T�[95|ZUEV�ZUEC\ZUFR�<JVCC��O<jV�IP,�CSC\�C�SGlJ�@I�9WE�B�:HTT�:R6l{L��CG{�IG[�oIPGS��RC,��DG�[H77�<6��:R85�JR66�JR7[R|R5-3{68|2�Z�@�Jml,|6|6\JR��\	P|4L�6�6u4��5�kNVDZ;R6+kR84<���4IP,�8��90���K�J9�\91��̫7X[KIP\JD0�F���CLI�lKCMS��J9��:STY,�T�O�:�@�K7�LNN.|ZORS<jJ��MZvZ|OLK�END�:uL�S��FVR�J�V3D,�KKPBV�\�APL�JAPV�ZCCG�:CCRvjCD�CDL̚wCSB�JCSK�j;CTK�CTB��\�D��\�C�z���CL�cTCLJ�l�TC��;TCZCTE�J���|�TE�J��<�TF*��F\�G��G��l�Hl�I�z)�l�k�C�TM\�M\�M��N*l�P,�P��R��;��TS��W��̚VGmF��P2��P2�z� �VPDFvLJVP;�VPR���VT�;� �JVTBZ��V�KIH�Vِ�M�<�VK,�V{�Gene�8�83EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W?�i?{?�7�0S�TD�4LANG�4�9�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~��������� �2�D�V�RBT�6OPTNm���� ����Ǐُ����!� 3�E�W�i�{�������ß�5DPN�4��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y��k�}ߏߡ߳�ted �4�8�������� 1�C�U�g�y���� ��������	��-�?� Q�c�u����������� ����);M_ q������� %7I[m �������/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ ����)�;�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ǯٯ������*�<�N�`�r����99���$FE�AT_ADD ?_	�������?  	��ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu������DEMO �Z��    ���}��'��0�]� T�f������������ ���#��,�Y�P�b� �������������� ��(�U�L�^����� �������ܯ��� $�Q�H�Z���~����� ���ؿ��� �M� D�Vσ�zόϦϰ��� �����
��I�@�R� �v߈ߢ߬������� ���E�<�N�{�r� ������������ �A�8�J�w�n����� ����������= 4Fsj|��� ���90B ofx����� ��/5/,/>/k/b/ t/�/�/�/�/�/�/�/ ?1?(?:?g?^?p?�? �?�?�?�?�?�? O-O $O6OcOZOlO�O�O�O �O�O�O�O�O)_ _2_ __V_h_�_�_�_�_�_ �_�_�_%oo.o[oRo do~o�o�o�o�o�o�o �o!*WN`z �������� �&�S�J�\�v����� �����ڏ���"� O�F�X�r�|������� ߟ֟����K�B� T�n�x�������ۯү ����G�>�P�j� t�������׿ο�� ��C�:�L�f�pϝ� �Ϧ�������	� �� ?�6�H�b�lߙߐߢ� ����������;�2� D�^�h�������� �����
�7�.�@�Z� d��������������� ��3*<V`� ������� /&8R\��� ������+/"/ 4/N/X/�/|/�/�/�/ �/�/�/�/'??0?J? T?�?x?�?�?�?�?�? �?�?#OO,OFOPO}O tO�O�O�O�O�O�O�O __(_B_L_y_p_�_ �_�_�_�_�_�_oo $o>oHouolo~o�o�o �o�o�o�o : Dqhz���� ���
��6�@�m� d�v�������ُЏ� ���2�<�i�`�r� ������՟̟ޟ�� �.�8�e�\�n����� ��ѯȯگ����*� 4�a�X�j�������Ϳ Ŀֿ����&�0�]� T�fϓϊϜ������� �����"�,�Y�P�b� �߆ߘ��߼������� ��(�U�L�^��� ����������� �� $�Q�H�Z���~����� ���������� M DV�z���� ���I@R v������ �//E/</N/{/r/ �/�/�/�/�/�/�/
? ?A?8?J?w?n?�?�? �?�?�?�?�?OO=O 4OFOsOjO|O�O�O�O �O�O�O__9_0_B_ o_f_x_�_�_�_�_�_ �_�_o5o,o>okobo to�o�o�o�o�o�o�o 1(:g^p� ������ �-� $�6�c�Z�l������� ϏƏ؏���)� �2� _�V�h�������˟ ԟ���%��.�[�R� d�������ǯ��Я� ��!��*�W�N�`��� ����ÿ��̿��� �&�S�J�\ωπϒ� �϶���������"� O�F�X߅�|ߎ߻߲� ���������K�B� T��x�������� �����G�>�P�}��t���������  ������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz�����y  �x�q� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p@������q�p�x���*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^��p���������������$FEAT_DEMOIN  ���� �����I�NDEX����ILECOMP [���B���8 SETUP2 \B�L�  N� w5_AP2B�CK 1]B	 � �)����%����E �	�� �5�Y�f� �B��x/�1/ C/�g/��/�/,/�/ P/�/t/�/?�/??�/ c?u??�?(?�?�?^? �?�?O)O�?MO�?qO  O~O�O6O�OZO�O_ �O%_�OI_[_�O__ �_�_D_�_h_�_�_
o 3o�_Wo�_{o�oo�o @o�o�ovo�o/A �oe�o���N �r���=��a� s����&���͏\�� �����"�K�ڏo��� ����4�ɟX������ #���G�Y��}�����0���ׯQ	� P�� 2� *.VRޯ(���*+�Q���0W�{�e��PC����>��FR6:��ؾg�����T   �2π���\� ��d�G*.F��ϕ�	óġ���o�ߓ�ST�M�9���ư%�d��ψߓ�HU߻�Jש�pf�x���GIF�A�L�-����ߑ��JPG����Lձ�n�����JS�H������6���%
JavaScriptt���CSe���Kֹ�v�� %Casca�ding Sty�le Sheet�s��j�
ARGN?AME.DT'��O�\;��[�k|�(k DISP* rUOп��� ��
TPEINS�.XML/�:\�CcCusto�m Toolba�r��	PASSW�ORD���FR�S:\�� %�Password Config/ c�Q/�J/�/���/:/ �/�/p/?�/)?;?�/ _?�/�??$?�?H?�? l?�?O�?7O�?[OmO �?�O O�O�OVO�OzO _�O�OE_�Oi_�Ob_ �_._�_R_�_�_�_o �_AoSo�_woo�o*o <o�o`o�o�o�o+�o O�os��8� �n��'���]� ����z���F�ۏj� �����5�ďY�k��� �����B�T��x�� ���C�ҟg������� ,���P��������� ?�ί�u����(��� Ͽ^�󿂿�)ϸ�M� ܿqσ�ϧ�6���Z� l�ߐ�%ߴ��[��� �ߣߵ�D���h��� ��3���W����ߍ� ��@����v���� /�A���e������*� ��N���r�����= ��6s�&�� \��'�K� o��4�X� ��#/�G/Y/�}/ /�/�/B/�/f/�/�/ �/1?�/U?�/N?�?? �?>?�?�?t?	O�?-O ?O�?cO�?�OO(O�O��F�$FILE_�DGBCK 1]����@��� < �)�
SUMMARY�.DG�OsLMD�:�O;_@Di�ag Summa�ry<_IJ
CONSLOG1__&Q_��_NQConso?le log�_HK	TPACCN�_�o%o?oJUTP� Account�in�_IJFR6�:IPKDMP.'ZIPsowH
�o�o�KU[`Except�ion�oyk'PME?MCHECK5o�_�*_K�QMemory DataL��F7l�)6qRIPE�_$6�Zs�%�q Pac�ket L�_�DL��$�	r�qSTA�T���S� �%�rStatuysT��	FTP�Ы�:���Vw�Qmment TBD؏�� >I)ETHERNE���
q��[�NQEthe�rn�p�Pfigu�ra�oODDCSVRF̏��ďݟd���� verif�y all��{D�{.���DIFF՟ໟ͟b��s��dif�fd��
q��CHG01Y�@�R��f�z�,��-?��2ݯį@֯k�v�����3a�8H�Z�� ������VTRNDIAG.LS�̿޿�s�^q3� Ope��q SQnost�icEW�)�VDEV7�DAT�t�Q�c�u�g�Vi�s��Device�Ϫ�IMG7ºo�����y��s�Ima�gߨ�UP��E�S��T�FRS:�\�� �OQUpd�ates Lis�t �IJg�FLEXEVENQ�X�j���f�F� UIF� Ev���B,��s�)
PSRB?WLD.CM��sL�������PPS_ROBOWEL���GLo�GRAPHICS4Dy�b�t����%4D G�raphics �Fileu��AO�;��rGIG����u�
YvGigE��ة�BN�? )}��HADOW������\sSha�dow Chan�g���vbQRCMERR�n��\s� CFG �Error�ta�il� MA���CMSGLIB ��"^o� �x��T�)��ZD����/Xw�ZD6 ad�HPNOTI���
/��/ZuNotif�ic��H/��AG UO�/yO?�O'?P?OO t??�?�?9?�?]?�? O�?(O�?LO^O�?�O O�O5O�O�OkO _�O $_6_�OZ_�O~_�__ �_C_�_�_y_o�_2o �_?oho�_�oo�o�o Qo�ouo
�o@�o dv�)�M� ����<�N��r� �����7�̏[���� ��&���J�ُW���� ��3�ȟڟi�����"� 4�ßX��|������ A�֯e�����0��� T�f����������O� �s��ϩ�>�Ϳb� �oϘ�'ϼ�K����� ��ߥ�:�L���p��� �ߦ�5���Y���}��� $��H���l�~��� 1�����g���� �2� ��V���z�	�����?� ��c���
��.��R d�����M� q�<�`� ��%�I�� /�8/J/�n/��/ !/�/�/W/�/{/?"? �/F?�/j?|??�?/?��?�?�$FILE�_FRSPRT � ���0�����8MDONLY 1]�5��0 
 �)�MD:_VDA�EXTP.ZZZ��?�?_OnK6%�NO Back? file 9O�4S�6Pe?�OOO�O �?�O__?>_�Ob_t_ _�_'_�_�_]_�_�_ o(o�_Lo�_po�_}o �o5o�oYo�o �o$ �oHZ�o~�� C�g��	�2�� V��z������?�ԏ��u�
���.�@��4VISBCKHA&C*.VDA������FR:\Z�ION\DATA\v�����Vision VD�B��ŏ ���'�5��Y��j� �����B�ׯ�x�� ��1���үg������� X���P��t���Ϫ� ?�οc�u�ϙ�(Ͻ� L�^��ς��)���M� ��q� ߂ߧ�6���Z� ����%��I��������:LUI_CONFIG ^�5�m��� $ 	h�F{�5�����`�)�;�I���|xq� s�����������a���  $6��Gl~ ���K���  2�Vhz�� �G���
//./ �R/d/v/�/�/�/C/ �/�/�/??*?�/N? `?r?�?�?�???�?�? �?OO&O�?JO\OnO �O�O)O�O�O�O�O�O _�O4_F_X_j_|_�_ %_�_�_�_�_�_o�_ 0oBoTofoxo�o!o�o �o�o�o�o�o,> Pbt���� ����(�:�L�^� p��������ʏ܏� ����$�6�H�Z�l�� ������Ɵ؟ꟁ��  �2�D�V�h������� ��¯ԯ�}�
��.� @�R�d����������� п�y���*�<�N� `����ϖϨϺ����� u���&�8�J���[� �ߒߤ߶���_����� �"�4�F���j�|�� �����[������� 0�B���f�x������� ��W�����,> ��bt����O���(:��  xFS�$�FLUI_DAT�A _���>��u�RESULT 2�`�� ��T�/wiza�rd/guide�d/steps/?Expertb� �//+/=/O/a/s/��/�/�*�Con�tinue wi�th G�ance�/�/�/??(?:?�L?^?p?�?�?�? �T-U��90� �� �?���9��ps�?0OBOTO fOxO�O�O�O�O�O�O �O� �_/_A_S_e_ w_�_�_�_�_�_�_�_�n�?�?�?�<Frip�Oo�o�o�o �o�o�o�o!3E _i{����� ����/�A�S�o�$on�HoAO�T�imeUS/DST[������+�=��O�a�s������'Enabl�/˟ݟ� ��%�7�I�[�m������T�?{�ݯ����Æ24Ώ3�E� W�i�{�������ÿտ 翦����/�A�S�e� wωϛϭϿ������π��Ưد� G��Region�χߙ� �߽���������)��;�+Americasou����� ��������)�;��?�y�#߅�G�Y��ditorL����� ��#5GYk}���+ Touch Panel ��� (recommen�)��� *<N`r��U��e�w��������accesd�./@/ R/d/v/�/�/�/�/�/��/Q|Conne�ct to Network�/(?:? L?^?p?�?�?�?�?�?(�?�?Y���������!/��Int?roducts߆O �O�O�O�O�O�O__ (_:_U^_p_�_�_�_ �_�_�_�_ oo$o6oHo e�Oeo?O� X_�o�o�o�o' 9K]o��R_� �����#�5�G� Y�k�}�����h`�ooj}oߏ�o��*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ 쯫���Ϗ1��X�j� |�������Ŀֿ��� ��0��A�f�xϊ� �Ϯ����������� ,�>���_�!���E��� ����������(�:� L�^�p���߸��� ���� ��$�6�H�Z� l�~���O߱�s����� �� 2DVhz ��������
 .@Rdv�� ������/��'/ ���`/r/�/�/�/�/ �/�/�/??&?8?� \?n?�?�?�?�?�?�? �?�?O"O4O�UO/ yO�OO?�O�O�O�O�O __0_B_T_f_x_�_ I?�_�_�_�_�_oo ,o>oPoboto�oEO�O iO�o�o�O(: L^p����� ��_ ��$�6�H�Z� l�~�������Ə؏�o �o�o�/��oV�h�z� ������ԟ���
� �.��R�d�v����� ����Я�����*� �������C����� ̿޿���&�8�J� \�nπ�?��϶����� �����"�4�F�X�j� |ߎ�M�_�q��ߕ��� ��0�B�T�f�x�� ������������ ,�>�P�b�t������� �������߱���%�� L^p����� �� $��5Z l~������ �/ /2/��S/w/ 9�/�/�/�/�/�/
? ?.?@?R?d?v?�?�/ �?�?�?�?�?OO*O <ONO`OrO�OC/�Og/ �O�/�O__&_8_J_ \_n_�_�_�_�_�_�_ �?�_o"o4oFoXojo |o�o�o�o�o�o�O�o �O�O�oTfx� �������� ,��_P�b�t������� ��Ώ�����(��o I�m��C�����ʟ ܟ� ��$�6�H�Z� l�~�=�����Ưد� ��� �2�D�V�h�z� 9���]���ѿ����
� �.�@�R�d�vψϚ� �Ͼ��Ϗ�����*� <�N�`�r߄ߖߨߺ� �ߋ�տ����#��J� \�n��������� �����"���F�X�j� |��������������� ������u7� ������ ,>Pbt3��� ����//(/:/ L/^/p/�/ASe�/ ��/ ??$?6?H?Z? l?~?�?�?�?�?��? �?O O2ODOVOhOzO �O�O�O�O�O�/�/�/ _�/@_R_d_v_�_�_ �_�_�_�_�_oo�? )oNo`oro�o�o�o�o �o�o�o&�OG 	_k-_����� ���"�4�F�X�j� |������ď֏��� ��0�B�T�f�x�7 ��[������� ,�>�P�b�t������� ��ί�����(�:� L�^�p���������ʿ ��뿭��џӿH�Z� l�~ϐϢϴ������� ��� �߯D�V�h�z� �ߞ߰���������
� �ۿ=���a�s�7ߚ� �����������*� <�N�`�r�1ߖ����� ������&8J \n-�w�Q���� ��"4FXj |�������� //0/B/T/f/x/�/ �/�/�/���/? �>?P?b?t?�?�?�? �?�?�?�?OO�:O LO^OpO�O�O�O�O�O �O�O __�/�/�/? i_+?�_�_�_�_�_�_ �_o o2oDoVoho'O �o�o�o�o�o�o�o
 .@Rdv5_G_ Y_�}_����*� <�N�`�r��������� yoޏ����&�8�J� \�n���������ȟ� ����4�F�X�j� |�������į֯��� �ˏ�B�T�f�x��� ������ҿ����� ٟ;���_�!��ϘϪ� ����������(�:� L�^�p߁ϔߦ߸��� ���� ��$�6�H�Z� l�+ύ�Oϱ�s����� ��� �2�D�V�h�z� ��������������
 .@Rdv�� ��}������� <N`r���� ���//��8/J/ \/n/�/�/�/�/�/�/ �/�/?�1?�U?g? +/�?�?�?�?�?�?�? OO0OBOTOfO%/�O �O�O�O�O�O�O__ ,_>_P_b_!?k?E?�_ �_{?�_�_oo(o:o Lo^opo�o�o�o�owO �o�o $6HZ l~���s_�_�_ ���_2�D�V�h�z� ������ԏ���
� �o.�@�R�d�v����� ����П������ ��]���������� ̯ޯ���&�8�J� \����������ȿڿ ����"�4�F�X�j� )�;�M���q������� ��0�B�T�f�xߊ� �߮�m��������� ,�>�P�b�t���� ��{ύϟ����(�:� L�^�p����������� ���� ��6HZ l~������ ���/��S�z �������
/ /./@/R/d/u�/�/ �/�/�/�/�/??*? <?N?`?�?C�?g �?�?�?OO&O8OJO \OnO�O�O�O�Ou/�O �O�O_"_4_F_X_j_ |_�_�_�_q?�_�?�_ �?�_0oBoTofoxo�o �o�o�o�o�o�o�O ,>Pbt��� ������_%��_ I�[���������ʏ ܏� ��$�6�H�Z� ~�������Ɵ؟� ��� �2�D�V��_� 9�����o�ԯ���
� �.�@�R�d�v����� ��k�п�����*� <�N�`�rτϖϨ�g� ����������&�8�J� \�n߀ߒߤ߶����� ���߽�"�4�F�X�j� |������������ ��������Q��x��� ������������ ,>P�t��� ����(: L^�/�A��e�� �� //$/6/H/Z/ l/~/�/�/a�/�/�/ �/? ?2?D?V?h?z? �?�?�?o���?� O.O@OROdOvO�O�O �O�O�O�O�O�/_*_ <_N_`_r_�_�_�_�_ �_�_�_o�?#o�?Go 	Ono�o�o�o�o�o�o �o�o"4FXio |������� ��0�B�T�ou�7o ��[o��ҏ����� ,�>�P�b�t������� iΟ�����(�:� L�^�p�������e�ǯ ��믭���$�6�H�Z� l�~�������ƿؿ� ���� �2�D�V�h�z� �Ϟϰ��������Ϸ� �ۯ=�O��v߈ߚ� �߾���������*� <�N��r����� ��������&�8�J� 	�S�-�w���c����� ����"4FXj |��_����� 0BTfx� �[��������/ ,/>/P/b/t/�/�/�/ �/�/�/�/�?(?:? L?^?p?�?�?�?�?�? �?�?����EO/ lO~O�O�O�O�O�O�O �O_ _2_D_?h_z_ �_�_�_�_�_�_�_
o o.o@oRoO#O5O�o YO�o�o�o�o* <N`r��U_� �����&�8�J� \�n�������couo�o 鏫o�"�4�F�X�j� |�������ğ֟蟧 ���0�B�T�f�x��� ������ү������ ُ;���b�t������� ��ο����(�:� L�]�pςϔϦϸ��� ���� ��$�6�H�� i�+���O��������� ��� �2�D�V�h�z� ���]���������
� �.�@�R�d�v����� Y߻�}����ߣ�* <N`r���� �����&8J \n������ ���/��1/C/j/ |/�/�/�/�/�/�/�/ ??0?B?f?x?�? �?�?�?�?�?�?OO ,O>O�G/!/kO�OW/ �O�O�O�O__(_:_ L_^_p_�_�_S?�_�_ �_�_ oo$o6oHoZo lo~o�oOO�OsO�o�o �O 2DVhz �������_
� �.�@�R�d�v����� ����Џ⏡o�o�o�o 9��o`�r��������� ̟ޟ���&�8�� \�n���������ȯگ ����"�4�F��� )���M���Ŀֿ��� ��0�B�T�f�xϊ� I������������� ,�>�P�b�t߆ߘ�W� i�{��ߟ���(�:� L�^�p������� ������$�6�H�Z� l�~������������� ����/��Vhz �������
 .@Qdv�� �����//*/ </��]/�/C�/�/ �/�/�/??&?8?J? \?n?�?�?Q�?�?�? �?�?O"O4OFOXOjO |O�OM/�Oq/�O�/�O __0_B_T_f_x_�_ �_�_�_�_�_�?oo ,o>oPoboto�o�o�o �o�o�o�O�O%7 �_^p����� �� ��$�6��_Z� l�~�������Ə؏� ��� �2��o;_� ��K��ԟ���
� �.�@�R�d�v���G� ����Я�����*� <�N�`�r���C���g� ��ۿ����&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲����ߕ��� ��˿-��T�f�x�� ������������� ,���P�b�t������� ��������(: ����A��� �� $6HZ l~=������ �/ /2/D/V/h/z/ �/K]o�/��/
? ?.?@?R?d?v?�?�? �?�?�?��?OO*O <ONO`OrO�O�O�O�O �O�O�/�O�/#_�/J_ \_n_�_�_�_�_�_�_ �_�_o"o4oE_Xojo |o�o�o�o�o�o�o�o 0�OQ_u7_ �������� ,�>�P�b�t���Eo�� ��Ώ�����(�:� L�^�p���A��eǟ ��� ��$�6�H�Z� l�~�������Ưد�� ��� �2�D�V�h�z� ������¿Կ������ �+��R�d�vψϚ� �Ͼ���������*� �N�`�r߄ߖߨߺ� ��������&��/� 	�S�}�?Ϥ������ �����"�4�F�X�j� |�;ߠ����������� 0BTfx7� ��[����� ,>Pbt��� �����//(/:/ L/^/p/�/�/�/�/�/ ����!?�H?Z? l?~?�?�?�?�?�?�? �?O O�DOVOhOzO �O�O�O�O�O�O�O
_ _._�/�/?s_5?�_ �_�_�_�_�_oo*o <oNo`oro1O�o�o�o �o�o�o&8J \n�?_Q_c_��_ ���"�4�F�X�j� |�������ď�oՏ�� ��0�B�T�f�x��� ������ҟ��� �>�P�b�t������� ��ί����(�9� L�^�p���������ʿ ܿ� ��$��E�� i�+��Ϣϴ������� ��� �2�D�V�h�z� 9��߰���������
� �.�@�R�d�v�5ϗ� Yϻ�}������*� <�N�`�r��������� ������&8J \n������� �����FXj |������� //��B/T/f/x/�/ �/�/�/�/�/�/?? �#�G?q?3�?�? �?�?�?�?OO(O:O LO^OpO//�O�O�O�O �O�O __$_6_H_Z_ l_+?u?O?�_�_�?�_ �_o o2oDoVohozo �o�o�o�o�O�o�o
 .@Rdv�� ��}_�_�_�_��_ <�N�`�r��������� ̏ޏ�����o8�J� \�n���������ȟڟ ����"����g� )�������į֯��� ��0�B�T�f�%��� ������ҿ����� ,�>�P�b�t�3�E�W� ��{�������(�:� L�^�p߂ߔߦ߸�w� ���� ��$�6�H�Z� l�~��������� �����2�D�V�h�z� ��������������
 -�@Rdv�� ������� 9��]����� ���//&/8/J/ \/n/-�/�/�/�/�/ �/�/?"?4?F?X?j? )�?M�?qs?�?�? OO0OBOTOfOxO�O �O�O�O/�O�O__ ,_>_P_b_t_�_�_�_ �_{?�_�?oo�O:o Lo^opo�o�o�o�o�o �o�o �O6HZ l~������ ���_o�_;�e�'o ������ԏ���
� �.�@�R�d�#���� ����П�����*� <�N�`��i�C����� y�ޯ���&�8�J� \�n���������u�ڿ ����"�4�F�X�j� |ώϠϲ�q������� 	�˯0�B�T�f�xߊ� �߮����������ǿ ,�>�P�b�t���� �������������� ��[�߂��������� ���� $6HZ �~������ � 2DVh'� 9�K��o����
/ /./@/R/d/v/�/�/ �/k�/�/�/??*? <?N?`?r?�?�?�?�? y�?��?�&O8OJO \OnO�O�O�O�O�O�O �O�O_!O4_F_X_j_ |_�_�_�_�_�_�_�_ o�?-o�?QoOxo�o �o�o�o�o�o�o ,>Pb!_��� ������(�:� L�^�o�Ao��eog� ܏� ��$�6�H�Z� l�~�������s؟� ��� �2�D�V�h�z� ������o�ѯ����� ˟.�@�R�d�v����� ����п����ş*� <�N�`�rτϖϨϺ� �����������/� Y���ߒߤ߶����� �����"�4�F�X�� |������������ ��0�B�T��]�7� ����m������� ,>Pbt��� i����(: L^p���e�w� �������$/6/H/Z/ l/~/�/�/�/�/�/�/ �/� ?2?D?V?h?z? �?�?�?�?�?�?�?
O ���OO/vO�O�O �O�O�O�O�O__*_ <_N_?r_�_�_�_�_ �_�_�_oo&o8oJo \oO-O?O�ocO�o�o �o�o"4FXj |��__���� ��0�B�T�f�x��� ����moϏ�o�o� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ���!��E�� l�~�������ƿؿ� ��� �2�D�V��z� �Ϟϰ���������
� �.�@�R��s�5��� Y�[���������*� <�N�`�r����g� ��������&�8�J� \�n�������c����� ������"4FXj |������� ��0BTfx� ���������� ��#/M/t/�/�/�/ �/�/�/�/??(?:? L?p?�?�?�?�?�? �?�? OO$O6OHO/ Q/+/uO�Oa/�O�O�O �O_ _2_D_V_h_z_ �_�_]?�_�_�_�_
o o.o@oRodovo�o�o YOkO}O�O�o�O* <N`r���� ����_�&�8�J� \�n���������ȏڏ ����o�o�oC�j� |�������ğ֟��� ��0�B��f�x��� ������ү����� ,�>�P��!�3�������$FMR2_G�RP 1a���� �C�4  B�[�	 �[�߿�ܰE��� F@ �5W�S�ܰJ���NJk�I'P�KHu��IP��sF!���?��  W�S�ܰ9��<9�8�96C'6<�,5���A��  �Ϲ�BHٳB�հ����@�33.�33S�۴߼�ܰ@UUT'�@���8��W�>u.��>*��<�����=[�B=����=|	<�K��<�q�=��mo���8�x�	7H<8�^�6�Hc7��x?����������"���F�X���_CFG� b»T �Q����X�NO {º
F0��� ��W�RM_CHKTYP  ���[�ʰ̰����ROM��_MIN�[����9����X��S�SBh�c�� ݶf�[�]������^�TP_DEWF_O�[�ʳ>��IRCOM����$GENOVR/D_DO.�d����THR.� dd���_ENB�� ^��RAVC��dO��Z� ���Fs�  G!� G����I�C�I(?i J���+��ĳ%����� ��QOU��j¼�������< 6�i�C�;]�[�?C�  D�+���@���B�����.��R SM�T��k_	ΰ\���$HOSTCh�19l¹[��d�۰� MC[����/Z�  27.�0� 1�/  e �/??'?9?G:�/j?�|?�?�?�,Z?T3	anonymouy  �?�?	OO-O?N�/ڰRHRK�/�?�O�/�O �O�O�O_V?3_E_W_ i_�O&_�?�_�_�_�_ �_@O�_dOvOSo�_�O jo�o�o�o�o_�o +=`o�_�_�� ���o&o8oJoL 9��o]�o��������o ɏۏ����4�j+� Y�k�}�������� � ��T�1�C�U�g� ����������ӯ��x� >��-�?�Q�c����� Ο���Ͽ���� )�;ς�_�qσϕϧ� ʿ ������%�7� ~�����߶ϣ���� �������Ϻ�3�E�W� i�ߍ��ϱ������� ��@�R�d�v�x�J��� ������������� +=`��������:$h!ENT� 1m P!\V  7  ?.c&�J�n ���/�)/�M/ /q/4/�/X/j/�/�/ �/�/?�/7?�/?m? 0?�?T?�?x?�?�?�? O�?3O�?WOO{O>O �ObO�O�O�O�O�O_ �OA__e_(_:_�_^_�_�_�_�ZQUICC0�_�_�_?odA1@oo.o�od2�o�lo~o�o!ROU�TER�o�o�o/!?PCJOG0�!192.168.0.10	o~�SCAMPRT�\!pu1yp��v�RT�o��� !�Softwar�e Operat�or Panel��mn��NAME� !�
!RO�BO�v�S_CF�G 1l�	 ��Auto�-started^'�FTP2�� I�K2��V�h�z��� ����ԟ����	� ��@�R�d�v���	��� ����:���)�;� M�_�&���������˿ �p���%�7�I�[� �"�4�F�ڿ����� ���!�3���W�i�{� �ߟ���D�������� �/�vψϚ�w�ߛ� �Ͽ���������+� =�O�a���������� ������8�J�\�n�p� ]�������� ��#5X�k }����0 /D1/xU/g/y/�/ RH/�/�/�/�//? �/??Q?c?u?�?�� �/?�?:/O)O;O MO_O&?�O�O�O�O�O �?pO__%_7_I_[_ �?�?�?t_�O�_O�_ �_o!o3o�OWoio{o �o�_�oDo�o�o�o�����_ERR �n��-=vPDU�SIZ  �`^��P�Tt>muWR�D ?΅�Q� � guest�f�������~�SCDMNG�RP 2o΅Wp��Q�`����fKL� 	P0�1.05 8�Q �  �|���  ;|��  �z[ ����w���*����>��x����[�ݏȏ��בP�Ԡ������)�����D�r���ت�p"�Pl�P���Dx��dx�*�����%�__GROU7�pLyN��	/�o����QUP��UTu�� �TYàL}�?pTTP_AUT�H 1qL{ <�!iPenda�n����o֢!KAREL:*������KC��ɯۯ���VISION SET�9���� P�>�h��f�������@���ҿ����X�CTRL rL}�O�uſa
��f?FFF9E3-ϝT�FRS:DEF�AULT��F�ANUC Web Server�� ��t�X���t@����1�C�U�g�;tWR_�CONFIG �s;� ��=qI�DL_CPU_P5C���aBȠP��w BH��MIN����q��GNR_IO�Fq{r�`Rx��NPT_SIM_DO���STAL_S�CRN� �.�I�NTPMODNT�OLQ����RTY�0����-�\�ENB�Q�-���OLNK 1tL{�p�������)�;�M���MA�STE�%���SL?AVE uL|��RAMCACHE�k�c�O^�O_CF1G������UOC���~��CMT_OP��8�PzYCL�������_ASG 1v;��q
 O�r� �������&8J\W�ENU�MzsPy
��IP�����RTRY_C�N��M�=�zs���bTu ������w���p/�p��P_ME�MBERS 2x�;�l� $��X"���?�Q'W/i)��RC�A_ACC 2y��  X�g� ��� 6��"�����&�#�#�/�����,�$BUF0�01 2z�= �fzu0  uW0f�:4�:4�:4U�:4�:4�:4�:3kgr4r4+a��oa�c,:3c<�4UM�4]�4o�4��4U��4��4��4Ò4iҒ4i4cq4d�4U�4&�46�4H�4UW�4i�4x�4��4U��4��4��4��4���4��4�:3e�rD rD0rDBrDS�rDerDurD�rD��rD�rDQDe�rDݪrD�:4:4:4$�:45:4G:4!Dfj:392$?63:1@1ER I0ERQ0ERY0ERa0ER i0ERq0:1x1}R�0}R�0Q �2:1�1�R �0�R�0�R�0�R�0�R �0�R�0�R�0�R�0�R �0�RrT�1:1�1�R@ �R	@�R@�R@�R!@ �R)@�R1@�R9@�RA@ �RI@�RQ@�RY@�Ra@ �Ri@�Rq@:1xA}b�@ }b�@}b�@}b�@}b�@ }b�@}b�@}b�@}b�@ }bZd�A}b�@}b�@ER �@ER�@ER�@ERPER@	PER*dQ:193-_ 65GSNrI2WSNrY2gS Nri2wS��x3�S�r�2 �P�2�S�r�2�S�r�2 �S�r�2�S�r�2�S�r �2�S�r�t�3c��	B c��B'c��)B7c�� 9BGc��IBWc��YBgc ��iBwc��xC�c���B �c���B�c���B�c�� �B�c��c��C�c���B �cNr�B�cNrRsNr�3�S'v��2{�4(r�}ŋ���<����po�o��2�HIS!2�}� ܷ! �2024-06-26����П���S  8�o�X
�`��;�Ql�)�;�M�_�o�/X�j���5�������Ư�� 7 h���h�j�����0�B�y��cN��1O��������� �_ 9 �cP��	�� ��$���mv��0��Y�k�}������Z�M 9 ,����mv��;M �� ������r��!Q�>� P�b�t߆ߘߪ߼��� ���)��(�:�L�^� p����������  ��$�6�H�Z�l�~� ��s��,P����K�������o�d�1�ޱd� 1_q� q���������ޱc�:��b>��A �A�CUgU�g��p���.  a>ٰ-/$/6/�H/6���~/�/�/��&�0@�A��;c"��o�c�/�/? ?����,?g?y?�?�? �?�?�?�?�?.?@?R? ?OQOcOuO�O�O�O�O �O�OO*O_)_;_M_ __q_�_�_�_�_��5p�����p/o$o6o�� �Td�VbF Vbro�o �o�o��o�o�Wd2r�2r��Vb �nocu�u��o �����B��B��qٰ�*�<�N�`� N/`/�����̏�Xc@����k�������Տ �.�@��O�O������ ����П�����*� a�s�`�r��������� ̯ޯ��9�K�8�J� \�n���������ȿڿ��ZI_CFG 2�~�[ H
C�ycle Tim}e�Busy��Idl��m�in�S�U�p��Read>(�DowG�C�����Cou�nt�	Num D�����̔���ީ�PROG����U�P�)/s�oftpart/�genlink?�current=�menupage,1133,1��C�U�g�y�Tä�SD�T_ISOLC ; �Y� ����J23_DSP_?ENB  ��T�~��INC ��������A   ?��  =���<#��
���:�o �2�D/�l���+OB��C��O������G_GROUP� 1���9<�*�����t�?"������Q'�L� ^�p�/�����������\�~�G_IN_�AUTO����PO�SRE���KANJI_MASK0���DRELMONG ��[�ϔ�y�� ������f��%����Ӕ�-���KCL_L N�UM��G$KEYLOGGINGD��P�!����LAN�GUAGE ��U��DE?FAULT ��Q�LG�����S�Ux� �8T�oH  ���'0������!�K͔�;���
*!(UT13:\ J/ L/Y/ k/}/�/�/�/�/�/�/��/$>(�H?�VLN�_DISP ����P�&�$�^4OCTOL0tDz����
���1GBOOK ��d4V�11�0�%O!O3OEOWO�iKyM�TËIgF	 �5)����O}���2�_BUFF 2�N�� ���2O� _�2��6_M�R_d_�_ �_�_�_�_�_�_�_o 3o*o<oNo`o�o�o�o��o���ADCS ������L�O���+=Oa�dIO ;2��k +��������� ���*�:�L�^�r� ��������ʏ܏����$�6�J�uuER_ITM��d������ ǟٟ����!�3�E� W�i�{�������ïկ������7x�SEVtD��t�TYP�ށ��s������)R�STe�eSCRN�_FL 2��}�����/�A�S�e�wϨ�TP{��b�}�=NGNAM�ԸE��dUPSf0G�I��2����_�LOAD��G �%��%DROP�_�EITO_3��ϑ�MAXUALcRMb2�@���9
K���_PR��2 � �3�AK�Ci0���qO=_'X�Ӭ�P �2��; �*V	Z����
* ��� 4��*��'�`�	xN� ��z��������� ��1�C�&�g�R���n� ����������	�� ?*cFX��� ����; 0q\����� ��/�/I/4/m/ X/�/�/�/�/�/�/�/ �/!??E?0?i?{?^? �?�?�?�?�?�?�?O OAOSO6OwObO�OD�wDBG*� ����ѢѤO�@_LDX�DISA����ssM�EMO_AP��E� ?��
  �A�H$_6_H_Z_l_~_��_�_K�FRQ_C_FG ����C�A �G@��S�@<��d%�\o�_�P��ݐ�����*Z`/\b **:eb�DXojho�F�o �o�o�o�o�o; �O��dZ�U�y|��z,(9�Mt�� �1��B�g�N���r� �������̏	����?�A�ISC 1���K` ��O�����O����O֟����K�]�_MSTR �3�~�SCD 1�]��l��{����� دïկ���2��V� A�z�e�������Կ�� �����@�+�=�v� aϚυϾϩ������� ��<�'�`�K߄�o� �ߓߥ��������&� �J�5�Z��k��� �����������F� 1�j�U���y������� ������0T?lx�MK�Q�,���Q�$MLTAR�M�R�?g�� ~s�@���@M�ETPU�@l���4�NDSP_A�DCOL�@!C�MNT7 *F�NSW(FSTLqIxi%� �,�����Q��*PO�SCF�bPR�PMV�ST51ݗ,� 4�R#�
g!|qg%w/�'c/�/ �/�/�/�/�/?�/? G?)?;?}?_?q?�?�?�?�?�1*SING_CHK  {�$MODA�S��e���#EDEV �	�J	MC:>WLHSIZE�Ml ��#ETASK �%�J%$1234?56789 �O�E�!GTRIG 1�,� l�Eo#_�y0_S_�}�FYP�A�u�9D"CEM_IN�F 1�?k`�)AT&FV0�E0X_�])�QE�0V1&A3&B�1&D2&S0&�C1S0=�])GATZ�_#o
dH'o Oo�QC_wohAo�o bo�o�o�o �_& �_�_�_o�3o��o ���o��"�4�� X���ASe֏ ���C�0���f� !���q�����s�䟗� ����͏>��b���s� ��K���w���ٯ� ɟ۟L����#����� Y�ʿ����$�߿ H�/�l�~�1���U�g� y����ϯ� �2�i�V� 	�z�5ߋ߰ߗ���PO�NITOR�G �?kK   	�EXEC1o�2*�3�4�5��@��7�8�9o ����(��4� ��@��L��X��d⠂�p��|��2��2���2��2��2��2���2��2��2��2*��3��3��3(�#A�R_GRP_SVw 1��[ (�1�@3>�?|�/��Q��6 `���@Q�>��z�RM�A_DsҔN��I_ON_DB-@�1M�l  �l s�FH"[+�l LFH��N BL"FI-ud1}E����)PL_NAM�E !�E� ��!Defaul�t Person�ality (from FD)b�*RR2�� 1��L�XL�p<�X  d�- ?Qcu���� ���//)/;/M/@_/q/�/�/�/f2) �/�/�/??,?>?P?b?t?f<�/�?�?�? �?�?�?
OO.O@OROHdOc	�6�?�N
�O�OfP�O�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_�O�O2oDo Vohozo�o�o�o�o�o �o�o
.@o!o v������� ��*�<�N�`�r���ޖ� F* GT?�G�Me���  �ÏՍfd �������(�6��� ���
 �m�~�h����� ������ğ֟ �����:���
�]�m�f��	`������|į��:�oAb	�����c A�  /���P���� r�������^�˿ݿȿ���%��R�� 1��	X ��, �� ��� a� �@D�  t�?��z�`�?f |�fA/���t�{	��;�	�l��	 ��xJ���x��� �� �<�@����� ��·�K��K ��K�=*�J���J���J9���
�ԏC߷�t��@{S�\��(E�hє��.��I���ڌ���T�;f�ґ�$��3���´  �@���>�Թ�$�  >̿���ӧUf�g�x`���� ��
���Ǌ��� _�  {x @T�}����  �H ��l�ϊ�-�	'�� � ��I� �  �<��+�:�È��È�=�����0Ӂ���N �[��n �@���f����f��k���,�av�  '������@2��@�0@�Ш����C��Cb C���\C������G��@������� )�Bb $/�!��L��Dz�o�ߓ�~��0��( �� -���������!����D�  ��恀?��ffG�*<� !}�q�1�8���B�>��bp��(�(���P��	������>�?����x����W�<
6b<���;܍�<����<���<�^���I/��A�{���fÌ�,�?fff�?_�?&� T�@��.�"�J<?�;\��"N\�3��� �!��(�|��/z��/j' ��[0??T???x?c? �?�?�?�?�?�?3��%F��?2O�?VO�/�wO�)IO�OEHG@� G@0��G�� G}ଙO�O�O_�	_B_-_f_Q_BL
��B[�Aw_[_�_b� �_�[�_��mO3o�OZo��_~o�o�o�o���bs��PV( @|po 	lo-*cU�ߡ!A���r5eCP�xLo�}?�����#��3��W�s���6�Cv�q�CH3� j�t����q������|^(hA� ��ALffA]���?�$�?���;�°u�æ��)�	ff��?C�#�
����g\)�"�33C��
�����<��؎G�B����L�B��s�����	";�H�ۚG���!G��WI�YE���C��+�8�I۪�I�5�HgM�G�3E��R�C�j=x�
�p�I���G��f�IV=�E<YD�C<�ݟȟ�� ��7�"�[�F��j��� ����ٯį���!�� E�0�i�T�f�����ÿ ���ҿ����A�,� e�Pω�tϭϘ��ϼ� �����+��O�:�s� ^߃ߩߔ��߸����� � �9�$�6�o�Z�� ~������������ 5� �Y�D�}�h����� ����������
C:.(䁳��/"����<��xt��q3�8��<��q4Mgu����q�VwQ�
4p�+4�]$ $dR�v���u%PD"P��Q�_/�Z/=/(/a/L+R�g/n/�/�/�/�/�/  %��/�/+??O? :?s?/�_�?�?�?�;�?�?O�? OFO4O�rLO^O�O�O�O��O�O�J  2 {FsH�GT�V�M�uBO�|r�pp�C��S@�R_�t@o}_�_f_�_�|\!�WɃ�_oo�(o�z?���@@*�z�D�p�pk1u�p�~
 6o �o�o�o�o�o�o );M_q�ڊsa� ����D���$MR_CAB�LE 2��� ]��T��LaMa?�PMaLb�p�%Z��&P�C�p�!�O4>�B���^�!Y4� �!�E�h\�&��v�_l  ��&P�v�^wdN�{0��$�s8ca��F��Q 6�H�XT��6Pv� C$�Č�]�n��	� 'z�g"������ �ɾ&P��C���=�u������� )z��~։��s 9��T�,�>���b��� ����Ɵ��Ο3�.�� P�(�:���^���j��#� �������pH�Z�l�*���** �sOM }��y���B�"��4�%% 23�45678901�ɿ۵ ƿ���� ��� AQ� �!
��z�not s�ent ���W��TESTF�ECSALG� e�g;jAQd��ga%�
,���@���$�r�̹������� 9�UD1:\mai�ntenance�s.xmS�.�@��vj�DEFA�ULT�\�rGRP� 2���  p�� �J�%  �%�1st mec�hanical �check��!����������E ��Z�(�:�L�^��"���controller�Ԍ��߰��D����� ��$�s�cM��L��""8b���v��B�����������/�C}�a�6����dv����s�C��ge��.� battery�&��E	S(:�L^p�	|�dui�z�ablet  �D�а�R����/"/4/s�>�greas��'f�r#-� |!�/�E��/�/�/�/�/s�
�oi,�g/y/�/�/t?�?�?�?�?"s��
�XֈW��1!<X�AO�E
c?8O JO\OnO�O�t��?O��'O�O_ _2_�D_s�Overh�auE��L��R !xXЌQ�_���O�_ �_�_�_oX�$�_0o����_o �_�o�o�o �o�oo�o?oQoco J\n���o� )��"�4�F�� �|��k��ď֏� ���[�0�B���f��� ��������ҟ!���E� W�,�{�P�b�t����� 矼����A��(� :�L�^�����ѯ㯸� �ܿ� ��$�s�H� ����~�Ϳ�ϴ����� ��9��]�o�Dߓ�h� zߌߞ߰�����#�5� G���.�@�R�d�v��� ������������� *�y���`���O���� ��������?�&u� J��n���� �);_4FX j|����% �//0/B/�f/� ��/��/�/�/�/? W/,?{/�/b?�/�?�? �?�?�??�?A?S?(O w?LO^OpO�O�O�?�O OO+O�O_$_6_H_ Z_�O~_�O�O�O�_�_��_�_o o�P�R	 T"oOoaoso�_�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ�x��
��  ��Q�?�  @�a �oW�i�{��fC������̟�h*�** �Q�V��� �2��D��h�z��������_�S������ կ7�I�[�����ɯ/� ��ǿٿ#���!�3� }�����{ύϟ��s� ������C�U�g��S� e�w�9ߛ߭߿�	����e�a�$MR_HIST 2��U}�� 
 \jR�$ 2345678901*�2����)�9c_���R�� a_���������=�O� a��*�x�����r��� ����9��]o &�J����� #�G�k}4���d�SKCFM�AP  �U������`���ONREL  ����лEXCFENB'q
��!FNC$/�$JOGOVLI�M'd�m �KE�Y'p%y%_P�AN(�"�"�RU�N`,p%�SF?SPDTYPD(%��SIGN/$TO1MOTb/!��_CE_GRP 1��U�"�:` ��n?�c[?�?�؆?�? ~?�?�?�?!O�?EO�? :O{O2O�O�OhO�O�O �O_�O/_�O(_e__ �_�_�_�_v_�_�_�_�o�׻QZ_ED�IT4��#TCO�M_CFG 1���'%to�o�o 
�Ua_ARC_!"���O)T_MN_M�ODE6�Lj_�SPL�o2&UAP�_CPL�o3$NO�CHECK ?^� � R dv������ ���*�<�N�`���NO_WAIT_�L 7Jg50NT]aѰ��UZ��_E�RR?12���ф ��	��-����R�d�ԍ��`O����| ��� 
aC w��Bb?�;Ӛ�8�t��,,N/A�@�W<� �� ?�j�ϟj�����قPARAMႳ.��N�
oQ�ph�o��� = e� ��������گ�ȯ���"�4��X�j�F�g�蜿��A�ҿ�"OD�RDSP�c6/(O�FFSET_CAqR@`�o�DIS���S_A�`ARK�7KiOPEN_FILE4�1�aKf�`�OPTION_I�O�/�!��M_PR�G %�%$*�����h�WOT��E7O����Z��  �  �Z"�÷"�	 �hW"�Z����RG_DSBL  ��ˊ���RIENTTO MZC���A(�z�U�`IM_D����O��V�LCT ���Gbԛa��Zd��_PEX��`7�*�RAT�g �d/%*��UP S���{��������������$PA�L�������_POS_CHU�7�����2>3�L�XLw�p��$� ÿU�g�y��������� ������	-?Q�cu����Y2 C���"4FX j|����� � //$/6/H/Z/l/~/�Y���.��/�/ςP�/??,?>? P?b?t?�?�?�?�?�? �?�?OO�/�/LO^O pO�O�O�O�O�O�O�O  __$_6_H_Z_)O;O �_�_�_�_�_�_�_o  o2oDoVohozo�o�o�_����o�m ���~BPw�m@�m���~�jw8� �w������2��T��p��w���H��t	�`���̏ޏ��:�o����� �2��pA�  I��j� `���������џ����@��#�)�O�r�1����� 8���,� �\Ԡ�� @oD�  ��?����~�?� ���!D�𕢒��%G�  ;��	l��	 �xJ젌������ �<:� ��� ��2��H(��H3k7�HSM5G�22�G���GN�3�%�R��oR�d�2�Cf��a��{�ׄ���������3��¸��4��>���К������3�A�q½{=q�!ª��ֱ� "�(«�=�2��� ��{  �@�Њ���  ��Њ�2��ς�	'� � ���I� �  ��V���=�������˖ß���  ��y��n @@"��]�<߭˄���䣟��N�Д�  '��Ь�w�ӰC��C��\C߰��Ϲ��߼�!���@�4��$�/��2�~�B��B� I�;�)�j客z+����쿱����������( �� -��#�������!��]�9��  q�?�ffaH�Z���C ��������8� �����>�|P��}�(� ��P�������^\�?��� x� ����<
6b<�߈;܍�<��ê<���<�#^�*�gv�A)ۙ��脣��F�?ff�f?}�?&� ��@��.��J<?w�\��N\��) ���������� �ޤy�N9r]� ������/&/ �J/5/n/�	g/��/c(G@ G@�0i�G�� G} ���/??<?'?`?K?\�?o?BLi�B��A�?y?�?|��?K�? ů�/QO�/xO�?�O�Ox�O�Om��b��n�t @|�O'_�OK_ 6_H_�_�3��A��RS�i�Cn_�_j_0O�]?��ooAo,o�ù�Wi���ToC���`CHQo>Jd�`a�a@I���>(hA� ��ALffA]��?�$�?����ź°u�æ��)�	ff���C�#�
�opg�\)��33C��
�����<���nG�B����L�B��s����	�0źH�ۚG���!G��WIY�E���C��+�½I۪I��5�HgMG��3E��RC��j=�~
�pI����G��fI�V=�E<YD�#Zo���
�� U�@�y�d��������� я�����?�*�c� N���r��������̟ ��)��9�_�J��� n�����˯���گ� %��I�4�m�X���|� ��ǿ���ֿ���3� �W�B�Tύ�xϱϜ� ��������	�/��S� >�w�bߛ߆߿ߪ߼� ������=�(�a�L�(q��)�y���Z����<���a3�8������a4Mgu�����aϴVwQ�(�4p?�+4�]B�B����p����������UPbP���QO%x�`1[FjR��������  C���I4mX��8
O������.//>/d/R/�Rj/|/�/�/�/�/��/:  2 F�s�gGT�&6�M�eBmp�R�P�aC��3@�_p?�?�? �?�?�?�=�S�O�O)O;OMO�c?��W�@@�j��`��`�1�`�^
 TO�O�O�O�O�O _#_5_G_Y_k_}_�_��_�j�A �����D��$PAR�AM_MENU �?B���  DE�FPULSE�[�	WAITTMO{UTkRCVo� SHELL�_WRK.$CU�R_STYL`�DlOPTZ1ZoP�TBooibC?oR_DECSN`���l �o�o�o&O J\n�������QSSREL_IOD  >�
1��u�USE_PROG %�Z%�@��sCCR` �
1�SS��_HOST !F�Z!X���M�T _���x������L�_TIMEb �h���PGDEBUG��p�[�sGINP_�FLMSK�E�T�� V�G�PGAr� 25��?��CHS�D��TYPE�\�0 ��
�3�.�@�R�{� v�����ï��Я�� ��*�S�N�`�r��� �������޿��+� &�8�J�s�nπϒϻ��G�WORD ?	��[
 	PR<2��MAI�`�gSU�a��TEԀ̒��	Sd�CO�L��C߸�L� UC�~�h�d*��TRACECTL� 1�B��Q� ��m n'���0�ށ�DT �Q�B��М�D� � ��qU���������1�@�@⨐��@�@� �� �	������Ҫ����&��.�Ӫ�������Ӫ&��.��6��>��*F�
H�H�H���u������� H� �����������������Ѫ����&��.��6��>�U�g�y���G������������ ���������� ��/�A�S�e�w�� �������������R������O��OAO�Ug�X��UXXXX�AXf����V�UV�V�V��V��UV��V��V��V���V��V�ѐ!�������@����  2DNhz�f� ���-�?����?�? �?����������d5(O :OLO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�N�`�r������� ��̏ޏ����&�8� J�\�n���������ȟ ڟ����"�4�F�P� $Or���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �f������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o��o�o�a�$PGT�RACELEN � �a  ����`��f_�UP ���e�q'pq p��a_CFG ��u	s�a p��LtLtfqwpqz�  �qu4rDEFSPD �?|��ap��`H_�CONFIG ��us �`j�`d�t��b �a��qP�t�q��`���`IN7pTRL ��?}_q8�u�P�E�u��w��qLt�qqv�`LID�8s�?}	v�LLB� 1��y 5��B�pB4Ńqv �އ؏	�s << �a?��'���A�o� U�w�������۟��ӟ@��#�	�+�Y�v�� ������ï
���������/�u�GRP 1�ƪ��a@��j��hs�aA��
D�� D@�� Cŀ @�٭^�t�q�����q�p���.� ���Ⱦ#´���ʻB�)��	���?�)�c��a>��>�,�������ζ� =49X=H�9��
���� @�+�d�O���s߬�o�x������  Dz���`
��8���H�n� Y��}��������� ����4��X�C�|����)��
V7.1�0beta1Xv� A�������!�����?!G��>\=y�#���{33A!���@��͵��8w�A��@� �A�s�@Ls���� ���"4FXLsAprLry�ā��_���@l��@�3�3q�`s��k���Anff�a���ھ��)�x�� �ar�T�n��t����	t�K�NOW_M  �|uGvz�SV ��z�r�&��� �>/�/G/�a���y�MM���{ ����	^u (�l+/�/',_t@7XLs����@���%�"4�.N�Vz�MRM��|-TU��y�c?u;eOAD?BANFWD~x�{STM�1 1�y��4Gar�ra_B�2Sem���?~s�;Co��2��O�7�3A�ntena_Full @��VOD e�qH��^OpO�O�O�O �O�O�O!_ __W_6_�H_�_l_~_�_�b�72��<�!4�_  �<�_�_N�3�_�_
oo�749oKo]ooo�7A5�o�o�o�o�76�o�o�772DVh�78�����7+MA�0��swwOVLD  �{��/a�2PARNUM  �;]��nu�SCH*� 8��
����ω�3�UP�D��[�ܵ+�wu_C�MP_r -��0�'��5C�ER_CHKQ����1�"e��N�`�RS>0�?G�_�MO�?_��#u__RES_G�0��{
Ϳ@�3�d�W��� {��������կ���@*�����P�� O��8`l�������` ��ʿϿ��`�	�� �1p)�H�M���ph� �ό���p��������V 1��5�1�!�@`y�ŒTHR_INR>0/�Z"�5�d:�MASSG� �Z[�MNF�y�MO�N_QUEUE ���5�6Ӑ~  *#tNH�U��N�ֲ؎��END�����EcXE�����BE��|����OPTIO�������PROGRAoM %��%���߰���TASK_�I,�>�OCFG �ά�]�����DAkTAu#�����Ӑ2�%B�T�f�x��� 5��������������,>P�INFO
u#� ������ ���'9K ]o���������/lx� � �;���ȀK_��q���S&ENB-�Hb-&q�&2�/�(G���2�b+ X,{		��=����/O��@��P4$�0���99)�N'_EDIT ���W?i?>��WERFL�-���3RGADJ ��F:A�  �5?@Ӑ�5Wј6��]!֐���?� ' Bz�WӐ<1Ӑ�%�%O�8;��50!�2��7�	H��l�0�,�BP�0��@�0�M*z�@/�B **:�B��O�F�O2��D��A �ЎO�@O	_,X��%�:��H�q��O$_@r_0_�_���Q@WA�� >]�_�_�_o�_o�_ �_
o�o.o�ojodovo �o�o�o�o�o�o\ XB<N�r�� ��4��0���&� ��J������������ �����x�"�t�^� X�j�䟎���ʟğ֟ P���L�6�0�B���f� ��������(�ү$�� ����>���z�t���  Ϫ������l�� h�R�L�^�DX	������0�� ���t$  :�L��o�
ߓߥ��7PREF ��:�0�0
�5IOR�ITYX�M6��1MPDSPV�:
B ��UT��C�6ODU[CT��F:��vNFOG[@_TG�0���J:?�HIBIT�_DO�8��TOE�NT 1�F; �(!AF_IN�E*�����!t�cp���!u�d��8�!ic�m'��N?�XY�3�vF<��1)� �A�����0������� ����' ]D �h������*>��3��9
BO8Tf�3>���2�B��G/�LC��4��;LFJAB,  ���F!//%/7/�5�F�Z�w/�/�/�/�3&ENHANCE �2
FBAH+d�?�%;�������Ӓ1�1PORT_NUM+���0���1_C_ARTRE�@��>q�SKSTA*��oSLGS�������C�Unothing?�?O�O�۶0TEMP ��N�"O�E�0_�a_seiban |߅OxߕO�O�O�O�O _�O'__K_6_H_�_ l_�_�_�_�_�_�_�_ #ooGo2okoVo�ozo �o�o�o�o�o�o1 U@e�v�� �������Q��<�u�.IVERSI�	�L��� d?isable�.GSAVE �N��	2670H7K71|�h��!�/0��9�:� 	^�4�$�ϐ����e��͟ߟ�����9�D�tC-Å_y� 1������ő�����Ǻ�URGE� B��r�WFϠ��-��9�W����l:W�RUP_DELA�Y �=n�WR_HOT %���7��/p��R_NORMALO�V�_�����SEMI���������QSKIPo��97��xf�=�b�a�s� ��H��ʹ��ø����� ���&��J�\�n�4� Fߤߒ������߲�� �� �F�X�j�0��|� �����������0� B�T��x�f�������|��ãRBTIF��5���CVTMOUڞ7�5���DC�Ro��� ��T�A�:CC��avC�>��;P>�[a:��_�H�� �c���^��?�S��`kϻ4��HϘ�� <
6�b<߈;܍��>u.�>*��<��ǪP0���2DVh z��������,GRDIO_TYPE  v��/�ED� T_CFGg ��-�BH]��EP)�2��+ ��B�u �/�* ��/�?�/%?=�/ V?�}?�Ϟ?���?�? �?�?�?O
O@O*Gl? qO��8O�O�O�O�O�O �O�O�O_<_^Oc_�O �__�_�_�_�_�_o �_&oH_Mol_o�oo �o�o�o�o�o�o�o" DoIho*j�� �����.3�E� �f� ���x������� �ҏ�*�/�N��b� P���t�����Ο��ޟ��:�+���R'INT� 2�R��!�1G;� i�{��"���8f�0 ��ӫ� �����M�;�q� W�������˿���տ �%��I�7�m��e� �ϑ��ϵ�������!� �E�3�i�{�aߟߍ� �߱���������A����EFPOS1 �1�!)  x���n#������� ������/��S��� w����6�����l��� ����=O����6 ���V�z�  9�]��� �Rd���#/� G/�k//h/�/</�/ `/�/�/??�/�/? g?R?�?&?�?J?�?n? �?	O�?-O�?QO�?uO �O"O4OnO�O�O�O�O _�O;_�O8_q__�_ 0_�_T_�_�_�_�_�_ 7o"o[o�_oo�o>o �o�oto�o�o!�oE W�o>���^ �����A��e�  ���$�����Z�l��� ��+�ƏO��s�� p���D�͟h�񟌟� '�ԟ�o�Z���.� ��R�ۯv�د���5� ЯY���}���*�<�v� ׿¿����Ϻ�C�޿�@�y��e�2 1� q��-�g�����	�� -���Q���N߇�"߫� F���j��ߎߠ߲��� M�8�q���0��T� ��������7���[� ����T�������t� ����!��W��{ �:�^p�� A�e �$ ��Z�~/�+/ ���$/�/p/�/D/ �/h/�/�/�/'?�/K? �/o?
?�?.?@?R?�? �?�?O�?5O�?YO�? VO�O*O�ONO�OrO�O �O�O�O�OU_@_y__ �_8_�_\_�_�_�_o �_?o�_co�_o"o\o �o�o�o|o�o)�o &_�o��B� fx��%��I�� m����,���Ǐb�� �����3�Ώ���,� ��x���L�՟p����� ��/�ʟS��w����<�ϓ�3 1��H� Z������6�<�Z��� ~��{���O�ؿs��� �� ϻ�Ϳ߿�z�e� ��9���]��ρ���� ��@���d��ψ�#�5� G߁�������*��� N���K����C��� g��������J�5� n�	���-���Q����� ����4��X�� Q���q�� �T�x� 7�[m�// >/�b/��/!/�/�/ W/�/{/?�/(?�/�/ �/!?�?m?�?A?�?e? �?�?�?$O�?HO�?lO O�O+O=OOO�O�O�O _�O2_�OV_�OS_�_ '_�_K_�_o_�_�_�_ �_�_Ro=ovoo�o5o �oYo�o�o�o�o< �o`�oY�� �y��&��#�\� ������?�ȏ����4 1�˯u����� ?�*�c�i���"���F� ���|����)�ğM� ����F�����˯f� ﯊�����I��m� ���,���P�b�t��� ���3�οW��{�� xϱ�L���p��ϔ�� �������w�bߛ�6� ��Z���~�����=� ��a��߅� �2�D�~� �������'���K��� H������@���d��� ��������G2k �*�N��� �1�U�N ���n��/� /Q/�u//�/4/�/ X/j/|/�/??;?�/ _?�/�??�?�?T?�? x?O�?%O�?�?�?O OjO�O>O�ObO�O�O �O!_�OE_�Oi__�_ (_:_L_�_�_�_o�_ /o�_So�_Po�o$o�o�Ho�olo�oۏ�5 1����o�o�olW ��o�O�s�� �2��V��z��'� 9�s�ԏ��������� @�ۏ=�v����5��� Y��}�����۟<�'� `��������C���ޯ y����&���J���� 	�C�����ȿc�쿇� ϫ��F��j�ώ� )ϲ�M�_�qϫ���� 0���T���x��u߮� I���m��ߑ����� ���t�_��3��W� ��{������:���^� ����/�A�{�����  ��$��H��E~ �=�a��� ��D/h�' �K���
/�./ �R/��/K/�/�/ �/k/�/�/?�/?N? �/r??�?1?�?U?g? y?�?O�?8O�?\O�? �OO}O�OQO�OuO�O�O"_t6 1� %�O�O_�_�_�_�O �_|_o�_o;o�__o �_�oo�oBoTofo�o �o%�oI�om j�>�b��� ����i�T���(� ��L�Տp�ҏ���/� ʏS��w��$�6�p� џ���������=�؟ :�s����2���V�߯ z�����د9�$�]��� �����@���ۿv��� ��#Ͼ�G�����@� �ό���`��τ�ߨ� 
�C���g�ߋ�&߯� J�\�nߨ�	���-��� Q���u��r��F��� j������������ q�\���0���T���x� ����7��[�� ,>x���� !�E�B{� :�^����� A/,/e/ /�/$/�/H/ �/�/~/?�/+?�/O?<5_GT7 1�R_�/ ?H?�?�?�?�/O�? 2O�?/OhOO�O'O�O KO�OoO�O�O�O.__ R_�Ov__�_5_�_�_ k_�_�_o�_<o�_�_ �_5o�o�o�oUo�oyo �o�o8�o\�o� �?Qc��� "��F��j��g��� ;�ď_�菃������ ˏ�f�Q���%���I� ҟm�ϟ���,�ǟP� �t��!�3�m�ί�� 򯍯���:�կ7�p� ���/���S�ܿw��� ��տ6�!�Z���~�� ��=ϟ���s��ϗ� � ��D������=ߞ߉� ��]��߁�
���@� ��d��߈�#��G�Y� k�����*���N��� r��o���C���g��� ��������nY �-�Q�u� �4�X�|b?t48 1�?);u ��/;/�_/� \/�/0/�/T/�/x/? �/�/�/�/[?F??? �?>?�?b?�?�?�?!O �?EO�?iOOO(ObO �O�O�O�O_�O/_�O ,_e_ _�_$_�_H_�_ l_~_�_�_+ooOo�_ soo�o2o�o�oho�o �o�o9�o�o�o2 �~�R�v�� �5��Y��}���� <�N�`��������� C�ޏg��d���8��� \�埀�	�����ȟ� c�N���"���F�ϯj� ̯���)�įM��q� ��0�j�˿��ￊ� Ϯ�7�ҿ4�m�ϑ� ,ϵ�P���tφϘ��� 3��W���{�ߟ�:� ����p��ߔ���A� ���� �:����Z� ��~�����=���a����� �����MA_SK 1����������XNO � ���� MOT�E  �R_C�FG �Y�����PL_RANG�UP���OWE/R ��� ��A��*SYST�EM*P�V9.3�044 �1/9�/2020 A� � ���RE�START_T �  , $F�LAG� $DS�B_SIGNAL�� $UP_C�ND4� �RS2�32r � �$COMMEN�T $DEVICEUSE4�PEEC$PAR�ITY4OPBI�TS4FLOWC�ONTRO3TI�MEOUe6CUz�M4AUXT���5INTERFA�CsTATU��  KCH� t $OLD�_yC_SW �'FREEFRO�MSIZ �AR�GET_DIR �	$UPDT�_MAP"� TS�K_ENB"EX�P:*#!jFAU�L EV!�RV�_DATA� � $n E� �  	$VALU�! 	j&GRP�_   �{!A  2 ��SCR	� �$ITP_�" $NUM� �OUP� �#TOT�_AX��#DSP��&JOGLI�F?INE_PCd��OND�%$U�M�K5 _MIR�1!4PP TN?8AsPL"G0_EXb0�<$�!� 814�!PG�w6BRKH�;&N�C� IS �  ��2TYP� �2�"P�+ Ds�#;0BSO�C�&R N�5DUM�MY164�"SV�_CODE_OP��SFSPD_O�VRD�2^LDlB3ORGTP; �LEFF�0<G� O�V5SFTJRUN�WC!SFpF5%3U�FRA�JTO�L�CHDLY7RE�COVD'� WS0* �0�E0RO��1�0_p@   �@��S NVER]T"OFS�@C� "FWD8A�D4A�1�ENABZ6�0TR�3$1_`1FDO>[6MB_CM�!FP=B� BL_M��!2hRnQ2xCV�"' �} �#PBGiW|8AM�z3\P��U�B�__MĀP�M� �1�AT$SCA� �PD�2�P�HBK+!:&aIOv�4 eIDX+bPPAj?a$iOd7e��U7a�CDVC_DBG"�a;!&�`�BD5�e1�j�S�e3�f^�@ATIO� ����AU�c� �S�A	B
0Y.#0�D�ȣX!� _�:&SU�BCPU%0SICN_RS�T, 1N|��S�T!�1$HW_C1�"]q.`�v�Q�$AT! � �$/UNIT�4�p�pATTRI= �r0�CYCL3NEC�A�bL3FLTR_2_FI9a7�c,�!LP;CHK_n�SCT>3F_�wcF_�|8��zFS+�R�rCHAGp�y�8�R�x�RSD�@'��1E#&7`_T�XP�RO�`@S�EMP'ER_0�3Tf�]p� f��P�DIA�G;%RAILAC4�c4rM� LO�0�A��65�"PS�"�2 X-`�e�SPR�`S. � �W�Ctaf	^�CFUNC�2�?RINS_T.!(0�w��� S_� �0��P�� 	d��WA�RL0bCBLCU	R��єAʛ�q͘Ƙ�DA�0���ѓʕL�D @,a3��!��8�3�TID�S��!� �$CE_RIA� !5AFDpPCX~��@��T2 �C9#̡b{QOI�pCVDF�_LE��#0(!�L�M�SFA�@HRD�YOL1	PRG8�H���>1(�ҥMUL�SE =#Sw3���$JJJ6BKGFKF�AN_ALMLV�3R�WRNY�HA#RD�0+&_P "��!2Q���!�5_�@:&�AU�Rk��TO_SBRvb��� ƺ�pvc�޳MPIN�F�@�q�)���REG'd~0V) 0R�C��1DAL_ \2F9L�u�2$MԐ(��#S��P� `�g�C�Mt`NF�qsONIP�qE�IPP� 9a$Y���!�"�!o� �o3EGP��#@��AR� �c�5�2�����|5AXE��'ROB�*RED&�&WR�@�1_=��3CSY�0ѥ0_�Si��WRI�@�ƅpST��#��0*@� �q	���3��� B� �A�ֺ3�D�POTO�� �@ARY�#��!���d�!1FI�0��$LINK��GT5H�B T_���A���6�"/�XYZt+"9�7G�OFF�@R�.�"���B� �l����A3$ ��F�I�p���4�4l��$_Jd�"(B�,a������8�"q����d��Ck6DUR���94�TURT�XZ�N����Xx��P��FL/�@s��l�P���30�"Q 1�� K
0M:$�53�]q7�SuD�Sw#ORQɆ�!�����Q7��0O[�ND�=#�!#�N1OVE8��M� ��R��R��Q!`P.!P! OAN}q 	�R����990� �b rJ9V����v��!ER1��	8�E��@n D�A��p��嘕Ă���v�AX�C�"��`�q�s ���0~3�~ F�~e�~�~E�~1��~Ҡ{Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�Ҡ��Ҡ�Ҡ�!)D7EBU}s$x���0삼!R*�AB�a�8A2V`|r 
 �"�c���%�Q7�7 �173�7F�7e�7 �7E�������LAB����yp�cGGRO�p��}��PB_ҁ ��̓��ð��6�1���5���6AND��8p�a3���-G �Q����AH�PH��p2�NTd��Cs@V�EL؁�}A��F��SERVEs@��� $����A!�!�@POR}�KP�иA� �B���	��]$�BTRQ�
�CdH��@
�G��2	�E�b��_  l8b��Q�ERR��R�I�P�@�FQTOQ�� L�}��YVĀ�G�E%�\ �DR}E�  ,�A��EP
�RA�Q �2 d�R7cܕU�@ ��$�F ׂ��m��CO�C��P  >8[COUNT�ђSFZN_CFG�AG 4�p%��rT\�zs�a�#`pJp�q�y�&c�� �� MGp+����`�OGp��eFAq����cX�8еk�ioQ��'ѴD�p8�Pz���HEL�A�-b 5���B_BAS\RSSR$�`�2�S�ѤL�!p1�W!p2Dz3�Dz4Dz5Dz6Dz7rDz8�WqROO��P�1�NL�� �AqB�C
�"pACK�&KIN�PT+�W�U��8	�k��y_PU8�~�|�OU�CP��%�s��Vl���YTPFWD_KARKQ-�:PRE�D�P����QUE$�Ā9 )���~���IU��#s/��8�@�/�SEM1ǆt1�A�aSTY�t3SO����DI�q��pQc��X��_TM9ßMANRQ �/�E�ND��$KEY?SWITCH2�G�����HE)�BEA�TMz�PE��LEPJR���0x�UF�F���G�S�DO_HOeM��Oz��pEF�PR��SbJі��uC⒐O��7P�QOV_�M��}�c�IOCM����1�BsHK��� D,�&�a`U�2R��M��a�r +�FwORC*�WAR���OM��  Q@�$�㰰U��P�Q1��g���3��4��T�@�POW�Lz��R�%�UNLO�0T��ED��  ��SNP��S.b �0N�ADDa`z��$SIZ*�$V�A�0�UMULTI�P�r���Az�? � $��Hƒ���SQc�1CFP�v�FRIFr�PS�w���ʔf�NF#�ODBUx�R@w������F��:�IAh�����������S"p�� g�  �cRTE��\�SGL.�T�x�&C`Gõ3a�/�S'TMT��`�P�����BW9 0�SHOW�h�qBANt�TP o���E������`mV_Gsb ��$PC�0�PoF�Bv�P��SP��A��p���@VD��rb�� �+QA002D.ҝ�6ק�6ױ��6׻�6�54�64�7�4�84�94�A4�B�4و�6ׇ17�}�6�F 4� ��@�����Z��T��t�1��1��1��U1��1��1��1��U1��1��1��23�U2@�2M�2Z�2g�U2t�2��2��2��U2��2��2��2��U2��2��2��33٨���M�3Z�3g�3�t�3��3��3��3���3��3��3��3���3��3��43�4�@�4M�4Z�4g�4�t�4��4��4��4���4��4��4��4���4��4��53�5�@�5M�5Z�5g�5�t�5��5��5��5���5��5��5��5���5��5��63�6�@�6M�6Z�6g�6�t�6��6��6��6���6��6��6��6���6��6��73�7�@�7M�7Z�7g�7�t�7��7��7��7���7��7��7��7���7��7���RVPzv�U�B �@��09r
�@V���A/ x �0R���+  �BM�@RP�`�4Q_�PR�@[U�A�R��DSMC��E�2F_U��=A��YS�L�P�@ �   �ֲ>g�������<iD��VALU>e�p�L�A�HFZAID_YL���EHI�JIh�?$FILE_ ��D��d$Ǔ�XCSA��Q h�0!PE_BLCKz�.RI�>7XD_CPUGY!� GY�Ic�O
TUB����R  � �PW`�p���QLA�n�S�Q�S�Q�TR?UN_FLG�U�T �Q�TJ��U�Q�T�Q�U�H��T`�T	 
w�T2L�_LIz��  �pG_�OT�P_ED�IU�_N/`�`7c� ?bة�pBQh�����TBC2 �! ��%�>��P��a�7aFqTτ�d݃TDC�PA�N`�`M�0�f�a&�gTH��U��d�3��gR�q�9�ERVAEЃt݃t	��a��p�` "X ;-$EqLENЃRt݃Ep�pRAv��Y@�W_AtS1Eq�D2&�wMO?Q�S���pI�.B�A�y�4Ep�{�DE�u��LACE� �CCC�.B��_�MA��v��w�T#CV�:��wT,�;� Z�P���s�~��sѕJ�A�M����JH���uā�uQq�2ѐ���݁�s�JK��VK�������	���J����JJv�JJ�AAL�@<��<�6��:�5�cm�N1a�m�,��D�L�p_\�Ű��ApC�F
�# `�0GRCOU�@J�Բ��N�`�C^�ȐREQUI9RrÀEBUu�Aqn��$T�p2"���Bp薋a	��d$ \�?@qhAPPR��C�LB
$H`N;�CLO}`K�S�e`��uv.`BCI�% �3��M�`�l��_M	G񱥠C �"P�����&���BRK��NO�LD����RTMO�6a�ޭ��J6`�P >��p��p��pZ��pc��p6+�7+�<�B��	@r�d&� ��lr��������PATH��������qxȪ����%0A��SCaAub��<���INDr�UC�p�q�C�U%M�Y�psP�����A q/ʤ�/�E�/�P�AYLOA�J2=L�0R_AN�apÁL�Pz�v�jɆ���R_F2LSHRt��LO{�R������>�ACRL_�qŐ����b�d�H�@B�$H��"�FLEX�>��aJ�f' P (��o�o+��>�Du( :Qcv�p ����fe��po��|F1���-������]�E��*� <�N�`�r�����4�Q� ������A�c���ɏۏ$���T��2�X:A�� �������� )�;�?�H�6�Z�c�u�p����>Ѭ�) ��``��˟ݟ�`�0ATF�𑢀EL��(a���J�(��JE۠C3TR��A�TN�1��HAND_VB�B>ѯ@�* $���F2���d�CS�W����+� $$M�����0ˡ�ڡ ������A�@g����A)��A���@˪A٫A� ��`P˪UD٫D�PȰG�P��)STͧ�!ک�!N�DY�P9����#% ��Fp���Ѫ���i����������P3�<�E�`N�W�`�i�r�MC�Ҏ�, ��ԓ� �n�5m��1ASYIMص.@�ض+A������_`��	�� �D�&�8�J�\�n�Ju�&��ʧC�I��S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R��&T ��3TWV�͢���&��ߪU��/�7�<ѓ`3HR`ta-��QLQ�1�DI��O�T8�b�P��. ; *"IAA*���$aG�2C�2cJ�$��I��P �/ � �MEB�� Mb�R4AT�PPT�@� ��ua���AP�l@zh�a�iT�@��� $DUM�MY1E�$PS�_D�RFॐ$��f3�FLA��Y�P���b}c$GLB_T��Uuu`1�p����EQa0 X(����ST����S�BR�PM21_V���T$SV_ERb��O_@KscsCLp�KrA��O'b�PGLv�@EW��1 4���a$Y|Z|W�s怯��AN`¼��qU�u2 ��N��p�@$GIU{}$�q 1u8�q�p��3 L���v�^B}$F^BE�vNWEAR��NK�F8����TANCK⥑JsOG��� 4`$JOINT�����uMSET��5�  �wE�H�� S������ ��6�k  MU��?���LOCK_FO�����PBGLVHG�L�TEST_X9M>���EMPt�[�q�r̀$U�Ќ�r��22���s,�3����Ҁ,�1MqCE����sM� $KAR���M�STPDRA8�pj�a�VEC��{��e�IU,�41�HE�ԀTOOL㠓Vv�RE��IS3��r��6N�A�ACH����5��O�}c�d3ڲ��pSI.� � @$RAIL_�BOXE��ppR�OBO��?�pqHOWWAR*���`�ROLM�bB����S��
�5���O_�F� !ppHTML5�Q����Щ�pڑ��7m� �R��O��8���v��z� �uOU��9 tpp(�14A��̀��PO֡%PIP��N��
�ڑ�S�,�����CORD�EDҀް̠5�XT<��q) �P� �O4` : D pOBP!"Ҁ{��j��cpj�^@$SYSj�ADR#�Pu`�TCH� ; M,��EN�RZ�Aف�_�t״��s�PV�WVAPa< �� p��r�UPRE�V_RT]1$E�DIT�VSHW�R�7v;���q��@D_`#R�+$HEADoA�Pl��A$�KE�q�`C�PSPD��JMP���L�UJ`R��dQ=r�O�϶I�S#�CiNE��$_T'ICK�AMX�\����HN-q> @pt������_GP֜�[�STYѲ�L�Oq�r��Ҩ�?j�
�Gݵ%$����t=7pS !$@Q��da�e!`�fP�0�SQUd� ��b�A�TERCy`Y��T=S�@ �pCp@����d�%Oz`�mcO�IZ�d�q�e�aPRM��a8����sPUQH�_DO=��ְXS��K�VAXiIg�f�1�UR� ���$#�Е��� _,����ET��Pۂ��J�5f�F�7g�A�!V�1�d9�2;� �SR|Al�о���#��5� �#��#�)#�)i� >'i�N'i�^&{����)�{����2��C����C`��WOiO{O�D���SCp B h�ppDS(�k��`SPL`�ATL �I����¼bADDRE�S��B'�SHIF���"�_2CH#r��I&p��TU&p�I� C��CU�STO��IaV��I�bDȲ,��0
��
�V�X�R`E \�����f�7���tC�#	���F���irt�TXSCR�EEl�F�P��T�INA�s�p��tp]����0G T�� fp,⧱eqBp&uᦲ8u�$#�RRO'0R��}�!�� 
	�;UE��H ��0��r�`S�q��RSMЂk�UV����V~!�PS_�s�&C�!�)�'C��Cǂz"� 2-G�UE�4Ibvr\�&8�GMTjPLDQ���Rp�z�	`BB�L_�W�`R`J ��f�>2O�qJ2L�E�U3"�T4RI;GH^3BRDxt�OCKGR�`�5TW�|�7�1WIDTH�H������a��� I�u�EY��QaK d��p��A�J�
�4�B�ACKH��b�5|q�X`FOD�GLAB�S�?(X`I�˂g$UR(�9@ �1�^`H4! L 8��QR�_k��\B_`R`�p͂����aACHB)O�R`M��w0�Uj0�CRۂM�LUqM�C��� ERV���p�0P<��4NV`��GE=B#���]�t��LP�E��E��Z)�Wj'Xz'XԐ&Y5*$[6$[7$[8	R��@�3�<���fԑŁ�S��M�1USR��tO <��^`U��r�rFO
�rP�RI��m����PT�RIP�m�U�NDO��P�p`��`m�4�l��#���� QWB�P7�G s�Tf�H�&RbOS�agfR��:">c��.qR��s�~�bH*�\!$�UQ.qS�o�o�#R)�>cOFFT���pT� �cOp� 1R�t/tS�GU��P.qx�Js�ETw�1SUB*� }f�E_EXE���V��>cWO>� eU�`^g��WA'���P�q!@� V_CDB�s�pݡ�PT�`�
�V�Q�r��OR���uRAU��tT��ͷ�q_���W 9|%�͸OWNA`޴$SRCE � ���D��\��MPFI8A�p��ESPD�� ����C���GƒG@+�5��!X `�`�r޴���COP�a	$��C`_w������rCT�3�q���qƲ� ���@� �Y"SHADOW��ઓ@�_UNSC�A��@��4M�DGD<ߑ��EGAC�,�ߡPG�Z (�0NO�@�D<�PE��B��VW�S�G|���![ � ���VEE#�aڒANG��$��c薴cڒLIM_X�c��c� � ���#��`� ��b�VF� �s�VCC�jв�\ՒC{�RA�lצ���RpNFA���%�E��Z2`G� ^0[�C`�DEĒ��� STE Q1���@�ꁻ@I��`�+0����`����P_A6�r���K��!]� 1Ҡ���A��\��сCPC�@�]�DRIܐ\�͑V�#Ѐ���D�TMY_UBY�T���c��F!���Y�븲����P_V�y��LN�B�MQ1$��DEY���EX�e��MUj��X�M� US�!���P_R��b�P� zߖG��PACIr� ʐf�ᔟ��c�´c��#�EqB��aWr8B����^ ܀�GΐP���\ C�R~``�_�0�@3!�1zri	�e�R�SW�� p�Yp��S�6�O�Q�1�A� X�#�E�UEd��Yp�pC�HKJ�`�@p���U� �EAN�ٖp�pXռ�`C�MRCV�!a� ��@O��M�pC«	��s����REF*7
��������/� �P��@���@��b�����_Y��ژ��ۣ�� Q$3������B��$b ����%���Q~��$GROU�  �c�����ʠ]��I�2^0��U` 0�_�I,�o � UL�ա`��C&�rAaB�?�NT�������� �A���Q��K�L����@õ��A���Q��T na$c t�`MD�p�8�HU���SA.�CMPE F  _�Rr�p@�����XS	 *�G�F/�b#d, &��@M�P^0۰UF_`C !���z �ROh0�"+���@���0C�UcREB���RI��
IN�p�����`d��d��ca�INE�H�y��0V�a-����3�W������0�C��i�LO�}��z�@0�!�QNSI ��݁���c$&�c$&.��X_PE-YW+Z�_M�ڒW�I��$�" �+R�'rRS�Lre �/�M�
`�RE�C7�G d�۰�̵ҭ�q���� u��Ȑ�������S_P�VnP ��I�A�vf �~pHD5R�p�pJO�P���$Z_UPz��a_LOW�5�1J�dA��LINubEP?�tc_i�1�1���@�G1@��V�x�g 5X�PA�THP X�CACH$�]E��yI�AT��{�C)�ID3FA�ETD�H��$HOD�pO�b@�{�d6��F�����p�PAGE�䁀VP�°�(RO_SIZ��2TZ3�`-X�0U�q�MPRZ���IMG���A9D�Y�MRE��R�7WGP��8�p��A�SYNBUF�V�RTD�U�T7Q�LE_2D-��U��`%CҡU1��Qu��U�ECCU��VEM��]EDb�GVIRC��Q�U�S�B�Q�LA|��p�NFOUN_�DIAG�YRE�X#YZ�cE�WѴh�8�dpqa`T��2�I�M�a�V|be��EGR�ABB��Y�a�LKERj�C4���FC-A�6504x��7u��S�BE��h'�`�CKLAS_@l�BA���N@i  G��T$��� @ݲմ$BAƠwj �!q�eb��uTYSp�H����2�šI�t:b�f��B)�E3VE����PK���flx��GI�pNO���2����qHO����k � ���
8��Pi�S�0ޗ��RO>�ACCEL?0=�-��VR_�U7@�`���2�p��AR��P�A��̎K�D��RE�M_But AB_�JMX �l�t�$SSC�U �"#�8��QN@m � ��S�P�NS� �VwLEX�vn T�ENAB 2�W@��oFLDRߨFI�P��t�ߨ(Ğ��2P}2HFo� ���V
Q MV_PI��8T@󐉰�F@�Z�+�#���8�8#��GA�B���LOO��J�CBx��w"SCON<(P�PLANۀ�Dp�3F�d�v�9PէAM��Q ;����SM0 E�ɥ�8ɥWb72�$`<�8T��,`RK<h"ǁVANC��@A�R_Ou N@p ( �-#<#c��c2���R_A/�N@q 4�������`	�^�
9
w�N@r hn��8�1^�&OFF`|�ap�`��`�DEA�Y
�P,`SK�DMP6�VIE��2q �w��@���rs < !{���4���r{7���D���
�CU�ST�U��t �$G�TIT1�$PR\��OPT<ap ��VSF�йsu�p�0`r&�*���MOwvI�|�ĄYJ�����eQ_WB��wI���� @O3��@�XVRxx�mr��T�� �Z�ABC��y �op����)�
�ZD�$�CSCH��z Lu����`�2�%PC ��7PGN ��<�<�A��_FUNH��@� 
�ZIPw�{I��LV,SL���~�� �ZMPCF��|��E����~X�DMY_LNH��=���M|��}� $�A� ]�CM+CM� C,SC&!���P�� $	J���DQ�������������_�Q,2�����UX�a\�UXEUL��a�������(�:�(�J���FTFqL��w��Z��~ *�6� �f���Y@Dp  8 $R�PyU��> EIGH��F��?(�iֱ��0��et� �a���F��$B�0�0@�	_SHIFD3-�ReVV`F�@��	$5��C�0��&!����D��b
�sx�uD��TR��V̱��Pr� H���!� ,���������4A�R�YP��%������%��   �%! � �H�(U N0���"�2������ɐ�q0GScPDak��� �P��O����0�ĬЯ�"!N�GVER`q �iw+I_A�IRPURGE { i  i/h�F`E�Tb� �+�  � h2ISO�LC  �,�"��!� �!�%��P+��_/*OB��Dm�?�@�!H?771  34n?��?�9� `�E/#�)x�� S232�� 1�i� L�TEk@ PEND�A�341 1D�3<*? M�aintenance Cons B��? F"O,DNo UseMJOO�nO�O�O�O�O2�2N�PO;/" 19%v�1CH=� �-�Q		9Q_!�UD1:___RS?MAVAIL/�/%��A!SR  ��+��H�_�P1�T7VAL.&���P�(.�YVL�}� 2|i�� D��P 	�/_oUQNo�o rci�o�g�o�o�o�o �o*,>tb �������� �:�(�^�L���p��� ����܏ʏ ��$�� H�6�X�~�l�����Ɵ ���؟�����D�2� h�V���z�������� ԯ
���.��R�@�b� d�v�����п����⿀��(�N�<�r�i��$SAF_DO_PULS. jQp�����CA� �/%��&0SCR ��`X���`�`
	14�1IAIE���b vo$�6�H�Z� l�~�ߢߴ������߬���HS��2�%�����d1�(�8�8rb��� @�"k� }���T�h� J`���_ @��T7 �����#�0�T D��0�Y�k� }��������������� 1CUgy�O<�Ef������  �5;�#o�� 1p�U��
�t��Di��������
  � ��*������gy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7O<A���`OrO�O�O�O�O �O�O�O?O�_._@_ R_d_v_�_�_�_�_�Q _�R0MJTo !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ JO��'�9�K�]�o� ������_ɟ۟��� �#�5�G�Y��_�U�_ �ҙ�����ϯ��� �)�;�M�_�m����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B�T�f�;�?�q߮� ����������,�>� P�b�t�������������������Y��	123456781�h!B!�)���F����� ������������  ��;M_q�� �����% 7I[l*��� ����//1/C/ U/g/y/�/�/�/n� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? O�/)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_O_�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�op_ �o�o�o/AS ew������ ���o+�=�O�a�s� ��������͏ߏ�� �'�9�K�]������ ����ɟ۟����#� 5�G�Y�k�}�������"��s�կ�w����0�L�CH  �Bpw�   ��=�2�� }� =�
���  	�o�ί���ǿٿ���r���� ��@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖ�%Ϻ��� ������&�8�J�\� n����������� ���"�Q�*������;�<M���D���  �]�w�*��Z򛱛�t  �d�����*�`*��$�SCR_GRP �1*P�3 � �*�� 6�	 �� 
��<�+*�'pUC|@��y�yD� W�!��y�	M-10�iA/7L 12�34567890ڙ�� 8��M1T� � �
�	L���	Č� N 
���Y���y�
M_	P������ ,��#H�
 ���1/�@A/g/y/H�ߙ! T/�/P/�/3��+���/B�S��,?*2C4r&Ad�R?  @0j5N?�7?��7&2R���?}:&F@ F�`�2�?�/�?�?O O-OSO>OwObO�O=�j1�2�O�O�O�O�DB��O�O;_&___J_�_ n_�_�_�_�_�_o�_ %o�5j�eSgxo6����uo�o�b�1�B̃|3�oh0�4j9j9B� w�$Y̯@HtA�Nhcu�/�%Ipp�drsq ����z�q�x� �.� (&�*�2� D�V�oz�e��������ECLVL  Ψ���iqpQ@���L_DEFAU�LT �����փHOT�STR�qq��MIPOWERF���H���WFDO�� �RVENT 1ɁɁ�� L!DUM�_EIP�����j�!AF_INEx‧���!FT}��֞����!-/� ���F�!RP?C_MAING�)�q�5���Y�VISb��t����ޯ!TP&ѠPUկ��dͯ*��!
PMON_POROXY+���e��v��D���fe�¿!�RDM_SRV�ÿ��g���!R�,*ϑ�h��Z�!
�[�M����iIϦ�!RLSYNC�����8����!R3OS|���4��>��!
CE�MTC�OM?ߓ�k-ߊ�!=	S�CONS�ߒ��ly���!S�WA'SRCݿ��m��"�;!S�USB#�n�n�!STMC��o]����� ѳ����,���P�V��ICE_KL ?�%d� (%S?VCPRG1S�����2�������o����4������5��6;@��7ch��H���9���� %��������0 ����X�����- ���U���}��� � /���H/���p/ ���/��F�/��n �/��?��8?�� �`?��/�?��6/�? ��^/�?��/X�j�� q���#OhO��lO�O{O �O�O�O�O�O�O _2_ _V_A_z_e_�_�_�_ �_�_�_�_oo@o+o doOo�o�o�o�o�o�o �o�o*<`K �o������ �&��J�5�n�Y����}���ȏ���^�_D�EV d���MC:�4����GRP 2�d���bx 	�� 
 ,V� ȡ�s�Z������� �����ߟ��@�'� 9�v�]�������Я��P��۫Y���� ܯI�1�4�]���j��� ��˿F�Ŀ��%�7� �[�B��f�xϵ�� !���A����ۿD�+� h�Oߌ�s߅��ߩ��� ��
���@�'�d�v��	y��^������ ����%��I�0�Y�� f�����8���������@��3��T7]�e �����)��
 �.@�dK�o@��!�9�� �!/G/���R/�/�/ �/�/�/"�/�/?? C?*?<?y?`?�?��? �?�?�?�?�?-OOQO 8OaO�OnO�O�O�O�O �O_�O)_;_"___�? �_�_L_�_�_�_�_�_ o�_7oo0omoTo�o xo�o�o�o�o�o! x_E�oU{b�� ������/�� S�:�w�^�p�����я��d �X�ZI�6 r��@�Z��0�+A�����dBj?BA�=��������B����AZ.�AĊ��+�A.�Q��B����5\���i6�A�u���'����%�Ꮛ�%PE�GA_BARRA�_ESTEIRA|����X�T����?=��=X���7
�?�>��A����������&���������Ax�P��f��U��'A�j������B�:��<�3����jB]+����T��%�T���d��ʐ���>�pc?���7�ԳT@�6��A�_���0n�����·�Ak���۸I�K9FA��G����B�!v,�-��C�3�����pBM�>�#�b�(�Y��������HX�?�L!���Q�B����AJ���Xk�@fD3���O�A��������Yw����.B�B��;��CH��z�B�?@���6���-Ϙ������n��=]����V@��?,������� վ��e�Ak�������OY�A������AB�J��;%�C$4�aƿBXZ9濠��
���ߘ�Ţ��� �ԭ(��^_���-\¯ԡ���گ���+����@��������ߔ�ᢧۙ�*נ�6��>�ԯb���zװ>
��BM��sﰲ�x�U<�߯�7@6|=���P�$�6��� N�@���b�G���L�}��������x7��~�K@���V��+A>r�r�F���������Y@+�@�<B���|�A�F�����B)���,o�?ɇ��~0��0~6��Z� Q�杚��������A�ߍ�]ܖA�?���������2[����>��ȥA��=�����NB ��$�w?�dj��to�7\�
`�.�%��Z�����A������*�@Ve�B� ������YN�#�B�D�	���9A����gB#
q�3���C4#��,??[BVM����COLOCA?_PRENS�����&//J/8/n/ \/~/�/�/�/�/ �/ ??D?2?T?�/�/ �?�/z?�?�?�?�?O 
O@O�?gO�?0O�O,O �O�O�O�O�O_ZO?_ ~O_r_`_�_�_�_�_ �_�_2_oV_�_Jo8o no\o�o�o�o�o
o�o .o�o"F4jX ��o��~�z� ��B�0�f����� V�����Џҏ��� >���e���.������� ��̟Ο���X�=�|� �p�^���������ȯ �D��T��H�6�l� Z���~�����ۿ��� Ϡ��D�2�h�Vό� ο���|�����
��� �@�.�dߦϋ���T� �߬���������<� ~�c��,����� �����D�)�;���� ��\������������ @���4"DFX �|����� �0@BT�� ��z��/�,/ /</���/�b/�/ �/�/�/?�/(?j/O? �/?�??�?�?�?�? �? OB?'Of?�?ZOHO ~OlO�O�O�O�OO�O >O�O2_ _V_D_z_h_ �_�_�O�__�_
o�_ .ooRo@ovo�_�o�o fo�obo�o�o* N�ou�o>��� ����&�hM�� ���n���������ȏ ��@�%�d��X�F�|� j��������,���<� ֟0��T�B�x�f��� ޟï��������,� �P�>�t�����گd� ο�����(��L� ��sϲ�<Ϧϔ��ϸ� ������$�f�Kߊ�� ~�lߢߐ��ߴ���,� �#�������D�z�h� ��������(��� 
�,�.�@�v�d����� �� �������( *<r�����b� ���$z� q�J����� �/R7/v /j/� z/�/�/�/�/�/*/? N/�/B?0?f?T?v?�? �?�??�?&?�?OO >O,ObOPOrO�O�?�O �?�O�O�O__:_(_ ^_�O�_�_N_p_J_�_ �_�_o o6ox_]o�_ &o�o~o�o�o�o�o�o Po5to�ohV� z����(�L �@�.�d�R���v��� ���$�����<� *�`�N���Ə���t� ޟp����8�&�\� ����L�����گȯ ����4�v�[���$� ��|�����ֿĿ�� N�3�r���f�Tϊ�x� �Ϝ����������� ��,�b�P߆�tߪ��� ��ߚ������(� ^�L���ߩ���r��� �� �����$�Z��� ����J����������� ��b���Y��2� z�����: ^�R�b�v� ���6�*// N/</^/�/r/�/��/ /�/?�/&??J?8? Z?�?�/�?�/p?�?�? �?�?"OOFO�?mOO 6OXO2O�O�O�O�O�O _`OE_�O_x_f_�_ �_�_�_�_�_8_o\_ �_Po>otobo�o�o�o �oo�o4o�o(L :p^��o�o� � ��$��H�6�l� ����\�ƏX�֏�� � ��D���k���4� ������ҟ���� ^�C����v�d����� ����ί��6��Z�� N�<�r�`��������� �󿪿̿���J�8� n�\ϒ�Կ�������� �������F�4�j߬� ����Z��߲������� ���B��i��2�� �����������J�p� A����t�b������� ����"�F���:�� Jp^������ � 6$Fl Z������� /�2/ /B/h/��/ �X/�/�/�/�/
?�/ .?p/U?g??@??�? �?�?�?�?OH?-Ol? �?`ONOpOrO�O�O�O �O O_DO�O8_&_\_ J_l_n_�_�_�O�__ �_o�_4o"oXoFoho �_�_�o�_�o�o�o �o0T�o{�oD �@�����,� nS�����t����� ����Ώ�F�+�j�� ^�L���p�������ܟ ��B�̟6�$�Z�H� ~�l����ɯۯ���� ����2� �V�D�z���������$SE�RV_MAIL + �����ʴ�OUTPUTո��@ʴRoV 2j�  㰧 (r����x��=�ʴSAVE����TOP10 2�� d 6 rƱ���϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t������n�YPY��FZN_CFG f��=��J���?GRP 2��g�� ,B   A� =�D;� B� �  B4=��RB21I�HELL��f�e�)��*�=�����%RSR����� �&J5G� k������.?�  ��/�>/P/"\/ ��X/z"{ �U'&"2��dh,g-�"EHKw 1S �/ �/�/�/#?L?G?Y?k? �?�?�?�?�?�?�?�?�$OO1OCO?OMM� S�ODFT?OV_ENBմ��e��"OW_REG�_UI�O�IMI_OFWDL~@�N��BWAIT�B �)��V��F�YwTIM�E��G_�VA԰_�A_UNcIT�C~Ve�LC�@WTRY�Ge�ʰ�MON_ALIA�S ?e�I%�he��oo&o8oFj�_ io{o�o�oJo�o�o�o �o�o/ASew "������� �+�=��N�s����� ��T�͏ߏ����� 9�K�]�o���,����� ɟ۟ퟘ��#�5�G� �k�}�������^�ׯ �����ʯC�U�g� y���6�����ӿ忐� ���-�?�Q���uχ� �ϫϽ�h������� )���M�_�q߃ߕ�@� �������ߚ��%�7� I�[�������� r������!�3���W� i�{���8��������� ����/ASe �����|� +=�as�� B����/�'/ 9/K/]/o//�/�/�/ �/�/�/�/?#?5?�/ F?k?}?�?�?L?�?�? �?�?O�?1OCOUOgO yO$O�O�O�O�O�O�O 	__-_?_�Oc_u_�_ �_�_V_�_�_�_oo�c�$SMON_�DEFPROG �&���Aa� &*S?YSTEM*obg� $JO0dR�ECALL ?}�Ai ( �}3�xcopy fr�a:\*.* v�irt:\tmp�back�a=>1�0.109.3.�21:11692� �a9228  a4bo�o�o	v}7�d�s:orderf?il.dat�l�o��odv�}.�bmgdb:�oA2 L���u2�e�o�o �d�a�s���q�o-� �oR�����,� P�a�s����3��N� ߟ�������L�]� o�����%�7�ʏ��� ���$���H�گk�}� ����=�ƟX�����  ���D�ֿg�yό��� /�¯T����ϊ��.� ����c�u߇ߚ�5߾� P������ϫϸ�N� _�q���'�9����������>��:pi�ckup_bar�ra_estei�ra.tp��em�p����[�m���<|�/�torno9���߉������5��lace��������d�v�};��sumir��6Q�Z�����",�prens 8���k}�"�1@CK�Z���=�furad/�U��e/w/
/���sem?_recep� 8/�J/�/�/�//#�co��/�/�/c?u?�? }�:��drop�"defeit�I?X?��?�?�8�:�4_1��?I�?hOzOOO_23OEOWO�O�O�O�O_3�O�O�Oh_z_� �1�D_U_�_�_�ߝ� �_���_dovo�o�� �Qo�o�o��o�o ���ofx�_�_�_= S���o�?o� b�t����o,9��o�� ������M^�p� ����0��ܟ� � �%���I�Z�l�~�����$SNPX_A�SG 2������� 7 0�%���Я�  ?���PAR�AM ��^�� �	��PӤ��Ө$�������OFT_KB_CFG  ӣ�����OPIN_S_IM  ����}���������RV�NORDY_DO�  )�U���QSTP_DSBi���ϐ�SR }�� � &#��D�O�O�:�TOP_ON_ERRʿ���o�PTN z�����A���RING_PRM�y�ܲVCNT_GOP 2��!���x 	�������#���Gߔ�VD��RP' 1��"�8Ѩ� *߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�}�z����� ����������
C @Rdv���� ��	*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?[?X?j?|?�? �?�?�?�?�?�?!OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLoso po�o�o�o�o�o�o�o  96HZl~ ��������� �2�D�V�`�PRG�_COUNTJ�9��{�ENB��}��M��L���_UPD� 1'�T  
k�����"�K�F� X�j���������۟֟ ���#��0�B�k�f� x���������ү���� ��C�>�P�b����� ����ӿο���� (�:�c�^�pςϫϦ� �������� ��;�6� H�Z߃�~ߐߢ����� ������ �2�[�V� h�z���������� ��
�3�.�@�R�{�v� ������������ *SN`r����t�_INFO {1�Ҁ� 	 ��3���)X@��>��L9 C� w�Bb?	��;ӛ8����,,MA�@�>�>�` AoB �@{w ?�� �>�@��a� ģ�C��Tp��1VC3�����"��3������YSD�EBUG��퀍d�Չ�SP_PAS�S��B?+LO�G ��� � � a�  ��с�UD1�:\;$�<"_MPACA-셽/�/�x!��/ 쁝&SAV D)��%d!|"�%��(SV�+TE�M_TIME 1�D'�� 0  z�#$ ��'�,5M7MEMBK'  �сd d/x�?�?�<X|Ҁg� @�?C�O :OJLOmOzI�J�%@p1�O�O�O�O "3 __$_6_H_Z_l_ �n_�_�_�_�_�_ �_�_o"o\�e1oVo hozo�o�o�o�o�o�o �o
.@Rdv0���O5SK�0�8����?���F1�� j�H2OJ�AJ�  @,4�A\O����(�O"�Oяb������p�O�  '� � ��0,:`� r���x_���3�Ο������$�C�7o g�y���������ӯ� ��	��-�?�Q�c�u�����������T1SVGUNSPD%%� '%��2M�ODE_LIM #a9"ܴ2�	�� D-۵ASK_?OPTION �9�!F�_DI ENB  �5%f��BC2_GRP 2!�u#o2��XB���C���ԼBCCF�G #��*< #6���`�@I� 4�Y��jߣߎ��߲� ��������E�0�i� T��x��������� ���/��S�>�w��� +�t���u�����c��� 	B-f�.��4 [ �������  02Dzh� ������/
/ @/./d/R/�/v/�/�/ �/�/�(���/?&?8? J?�/n?\?~?�?�?�? �?�?�?O�?4O"OXO FOhOjO|O�O�O�O�O �O�O__._T_B_x_ f_�_�_�_�_�_�_�_ oo>o�/Voho�o�o �o(o�o�o�o�o( :Lp^��� ����� �6�$� Z�H�~�l�������؏ Ə��� ��0�2�D� z�h���To��ȟ��� 
���.��>�d�R��� ����z�Я������ �(�*�<�r�`����� ����޿̿���8� &�\�Jπ�nϐϒϤ� �����ϴ��(�F�X� j��ώ�|ߞ��߲��� �����0��T�B�x� f������������ ��>�,�N�t�b��� �������������� :(^�v��� �H���$H Zl:�~��� ����2/ /V/D/ z/h/�/�/�/�/�/�/ �/?
?@?.?P?R?d? �?�?�?t�?�?OO *O�?NO<O^O�OrO�O �O�O�O�O�O__8_ &_H_J_\_�_�_�_�_ �_�_�_�_o4o"oXo Fo|ojo�o�o�o�o�o �o�o�?6Hfx ���������v&��$TBCS�G_GRP 2$��u� � �&� 
 ?�  Q�c�M���q� �������ˏ��*��1�&8�d, ��F�?&�	 HCwA����b�~�CS�B�I�x����V�>��ͪ��n�Ќ�ԝB��3�33��Blt�������AÐ�ff1f:��.�C���=�l�?����G�w�R���A&��̧�����@��I��-��� 
�X�u�@�R�����̻������	V3.�00I�	mt7���*� �%��ֶY��@ff&�5 &�H�� N� ��O�  ����Ͱ ϏϘ�*�J21�'�8��Ϥ�CFG [)�uB� E�V�����d���#��#�I�W��p W�}�hߡߌ��߰��� �����
�C�.�g�R� ��v��������	� ��-��Q�<�u�`�r� ����������I�cp "4��gRw� �����	- ?�cN�r�� &������/</ */`/N/�/r/�/�/�/ �/�/?�/&??J?8? Z?\?n?�?�?�?�?�? �?O�? OFO4OjOXO �O�O`�O�OtO�O_ �O0__T_B_x_f_�_ �_�_�_�_�_�_�_,o oPoboto�o@o�o�o �o�o�o�o�o(L :p^����� ��� �6�$�F�H� Z���~�����؏Ə�� ��2��OJ�\�n�� ������������ 
�@�R�d�v�4����� ����ί����ү(� N�<�r�`��������� ʿ̿޿��8�&�\� Jπ�nϐ϶Ϥ����� ����"��2�4�F�|� jߠߎ����߀��� � �߼�B�0�f�T��x� ������������ >�,�b�P��������� v�������:( ^L�p���� � �$H6l Z|������ /�/ /2/h/�߀/ �/�/N/�/�/�/
?�/ .??R?@?v?�?�?�? j?�?�?�?�?O*O<O NOOO�OrO�O�O�O �O�O�O _&__J_8_ n_\_�_�_�_�_�_�_ �_o�_4o"oXoFoho �o|o�o�o�o�o�o �/$6�/�oxf� �������,� >���t�b������� Ώ��򏬏��&�(� :�p�^���������ܟ ʟ�� �6�$�Z�H� ~�l�������دƯ�� � ��D�2�T�z�h� ��Jȿڿ������ 
�@�.�d�Rψ�vϬ� �����Ϡ������ *�`�r߄ߖ�Pߺߨ� ���������&�\� J��n�������� ����"��F�4�j�X� z�|����������� ��0B�Zl~( �������, Pbt�D��p����   �# &0/"��$TBJOP_G�RP 2*���  ?��&	H"O#,V,����� ��� =k%  Ȯ� � �� �$� @ g"	 ��CA��&��S�C��_%g!�"G;��"k��/�+�=�CS�??��?�&0%0?CR  B4�'??xJ7�/�/?333�2�Y&0}?�:;��v� 2�1�0-1*20��6?�?20��7C� � D�!�,� BL���OK:�Z��Bl  @pB@�^� s33C�1 �?�gO  A�zG�2�jG�&)A)E�O�J;���|A?�ff@,U@�1C�Z0zjO�O�z@���U�O�$f�ff0R)_;^;xCsQ?ٶ4)@�O�_�tF�X_J\EU�_�V:'�t-�Q(B�*@�O oh�&-h$oZGLo6o Doro�o~o8o�o�o�o �o3�oRlVPd��V4�&`�q��%	V3.00�m#mt7A@�s*��l$!�'� �E��qE����E�]\E�H�FP=F�{�F*HfF@D��FW�3Fp?�F�MF����F�MF���F�şF���F�=F����G�G.�8�CW�RD3l�)D��E"���Ex�
E���E�,)Fd�RFBFHFn�� F��F���MF�ɽF�,�
GlGg�!G)�G=���GS5�Gi���;��
;�Uo�|& : @XzQ&/��&"��?�0�&=;-ESTPARS  (�a E#HRw�ABL�E 1-V) $@�#R�7� � �
R�R�R�'#!R�	R�
R�R���!UR�R�R���'RDI��`!�� ԟ���
�r�Oz���@������̯ޮ��Sx�^# <�����ÿտ� ����/�A�S�e�w� �ϛϭϿ�������;- w�{�_"��6��1�C� U���%�7�I�[���~�NUM  ��`!� $  ���m���_CFG �.���!@H IMEBF_TT}�0��^#��G�VE10m��H�]�G�R 1/��� 8�"d �� �A�  �� ����������� �2� D�V�h�z��������� ����/
e@R hv������ �*<N`r ������'// /]/8/J/`/n/�/�/��/�/r���_��t�@�~�t�MI_CH�ANS� ~� !3D_BGLVLS�~��s�$0ETHERA�D ?��w0�"��/�/�?�?l�$0oROUTq�!��!�4�?�<SNM�ASKl8~�}1255.2E�s0OBOTO��st�OOLOFS�_DI}��%V9O�RQCTRL !0���#��MT�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo�&l�OIo8omoq�PE?_DETAIJ8�J�PGL_CONF�IG 6����/cell/�$CID$/grp1qo�o�o/壀�?Zl~�� �C���� �2� �V�h�z�������?� Q����
��.�@�Ϗ d�v���������M�� ����*�<�˟ݟr�@��������̯@�}a� ��&�8�J�\���^o��c��`���˿ݿ� ��Z�7�I�[�m�� �� ϵ���������� !߰�E�W�i�{ߍߟ� .������������ A�S�e�w����<� ��������+���O� a�s�������8����� ��'9��]o ����F��� #5�Yk}�����`�U�ser View� �i}}1234?567890�/ /,/>/P/X$� �cx/���2�U�/�/��/�/??s/�/�3 �/b?t?�?�?�?�??�?�.4Q?O(O:OLO ^OpO�?�O�.5O�O �O�O __$_�OE_�.6�O~_�_�_�_�_�_7_�_�.7m_2oDoVo@hozo�o�_�o�.8!o �o�o
.@�oa�gr lCamera��o�@���� �ޢE� *�<�N��h�z��������I  �v�)� �$�6�H�Z�l���� ������؟���� �2�Y��vP9ɟ~��� ����Ưد���� � k�D�V�h�z�����E� W�I5����� �2� D��h�zό�׿���� ������
߱�W�ދ�� X�j�|ߎߠ߲�Y��� ����E��0�B�T�f� x�߁ulY������� ��
����@�R�d��� ��������������W�  iy�.@Rdv� /����� *<N��W��i�� ������/*/ </�`/r/�/�/�/�/as9F/�/??1? C?U?�f?�?�?D/�?��?�?�?	OO-O�j	�u0�?hOzO�O�O�O �Oi?�O�O
_�?._@_ R_d_v_�_/OAO�p�{ ,_�_�_oo)o;o�O _oqo�o�_�o�o�o�o �o�_�u���oM_ q���No��� :�%�7�I�[�m� NEa����ˏݏ�� ��7�I�[������ ����ǟٟ����ͻp� %�7�I�[�m��&��� ��ǯ�����!�3� E�쟒�9�ܯ������ ǿٿ뿒��!�3�~� W�i�{ύϟϱ�X��� ��H����!�3�E�W� ��{ߍߟ����������������   ��L�^�p������������ ��   "�*�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/�r/�/�  
��(�  �@�( 	 �/�/�/�/�/?  ?6?$?F?H?Z?�?~?д?�?�?�*2� �l�O/OAO��eOwO �O�O�O�O��O�O�O _TO1_C_U_g_y_�_ �O�_�_�__�_	oo -o?oQo�_uo�o�o�_ �o�o�o�o^opo M_q�o���� ��6�%�7�~[� m���������ُ� ��D�!�3�E�W�i�{� ԏ��ß՟���� �/�A�S���w����� ⟿�ѯ�����`� =�O�a����������� Ϳ߿&�8��'�9π� ]�oρϓϥϷ����� ����F�#�5�G�Y�k� }��ϡ߳�������� ��1�C�ߜ�y�� ������������	�� b�?�Q�c�������� ������(�)p� M_q������0@ �������� ��#fr�h:\tpgl\�robots\m�10ia4_7l.xml�Xj| �������.��/1/C/U/g/y/ �/�/�/�/�/�/�// ?-???Q?c?u?�?�? �?�?�?�?�?
?O)O ;OMO_OqO�O�O�O�O �O�O�OO _%_7_I_ [_m__�_�_�_�_�_ �__�_!o3oEoWoio {o�o�o�o�o�o�o�_ �o/ASew� ������o�� +�=�O�a�s����������͏ߏ�I� �<<  ?��4�� ,�N�|�b�������ʟ �Ο���0��8�f� L�~���������������(�$TPG�L_OUTPUT� 9����� $�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}π�ϡϳ�����$�����2345678901��� �2�D� V�^����υߗߩ߻� ����w����'�9�K�]���}g������ ��o����1�C�U� g���u����������� }���-?Qc�� ������� );M_q	 �������%/ 7/I/[/m///�/�/ �/�/�/�/�/?3?E? W?i?{??%?�?�?�? �?�?O�?OAOSOeO wO�O!O�O�O�O�O�O�_�O� $$Ӣ��OW=_o_a_�_ �_�_�_�_�_�_�_#o oGo9oko]o�o�o�o �o�o�o�o�oC5g}��������}@��"�� ( 	 i W�E�{�i�����Ï�� ӏՏ���A�/�e� S���w��������џ ���+��;�=�O����s����Ƹ  <<\ޯ�)�ͯ �)��M�_���ʯ�� ��<���ؿ��Ŀ� � ~�$�V��BόϞ�x� ����2ϼ�
ߤ���@� R�,�v߈���p߾��� j�������<�߬� r��������� �`�&�8���$�n�H� Z�������������� "4Xj��R� �L����| Tf ��v� �0B//�&/P/ */</�/�/��/�/h/ �/??�/:?L?�/4? �??n?�?�?�?�? O ^?�?6OHO�?lO~OXO �O�OO$O�O�O�O_ 2___h_z_�O�_�_ J_�_�_�_�_o.o���)WGL1.X�ML�cm�$TP�OFF_LIM �Š�p����qfN_SVy`  ��t�jP_MOoN :���d��p�p2miSTRTCHK ;���f~tbVTCO�MPAT�h*q�fVWVAR <�m�Mx�d  �e�p�bua_D�EFPROG �%�i%COL�OCA_MESA_IRVISI�`��rISPLAY��`�n�rINST_�MSK  �| ��zINUSER� �tLCK)��{Q?UICKME�pO�ޕrSCREl����+rtpsc@�t)������b��_���STz�iRACE_CFG =�i�Mt�`	nt
?���HNL 2>�z���T{ zr@�R� d�v���������К�ITEM 2?,�� �%$1234567890�%�  =<�C�U�]�  !c�k�wp'���ns�ѯ5��� �k������j�ů�� 鯕���A�1�C�U�o� y�󿝿I�oρ�忥� 	��-ϧ�Q���#�5� ��A߽�����e߳�� ����M���q߃�L�� g��ߋ����%�w�  �[���+�Q�c��� o��������3��� {�;������G_ ����/�Se. �I�m�� �=�a/3/� �����k//�/ �/�/]/?�/�/�/? �/u?�?�??�?5?G? Y?�?+O�?OOaO�?mO �?�?�OO�OCO__ yO+_�O�Ox_�O�_�O �_�_�_?_�_c_u_�_ o�_Wo}o�o�_�oo )o;o�o�oqo1C�o O�o�o��%���[��Z��S��@��_��  ے_� ����y
 Ï�Џ����UD1:\����q�R_GRP �1A �� 	 @�pe�w�a��� ������ߟ͞�����ّ�>�)�b�M�?�  }���y����� ӯ������	��Q� ?�u�c���������Ϳ��	-���o�S�CB 2B{� h�e�wωϛϭϿ��������e�UTOR?IAL C{���@�j�V_CONFIG D{����������O�OUTPU�T E{�����������%�7� I�[�m������� ��������%�7�I� [�m������������ ����!3EWi {�������� /ASew� ������// +/=/O/a/s/�/�/�/ �/�/��/??'?9? K?]?o?�?�?�?�?�? �/�?�?O#O5OGOYO kO}O�O�O�O�O�O�? �O__1_C_U_g_y_ �_�_�_�_�_�O�_	o o-o?oQocouo�o�o �o�o�o�_�o) ;M_q���� ��yߋ����-�?� Q�c�u���������Ϗ ���o�)�;�M�_� q���������˟ݟ�  ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ���
��/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������� 1CUgy��� ����	-? Qcu��������/�x���$/6/ !/a/��/ �/�/�/�/�/�/?? '?9?K?]?�?�?�? �?�?�?�?�?O#O5O GOYOkO|?�O�O�O�O �O�O�O__1_C_U_ g_xO�_�_�_�_�_�_ �_	oo-o?oQocot_ �o�o�o�o�o�o�o );M_q�o� �������%� 7�I�[�m�~������ Ǐُ����!�3�E� W�i�z�������ß՟ �����/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿����'�9�K�]�o�~��$�TX_SCREE�N 1F8%;  �}�~��� ������
����m& ��\�n߀ߒߤ߶�-� ?������"�4�F�� j��ߎ��������� _����0�B�T�f�x� ������������ ��>��bt�� ��3�W( :L^����� ���e/�6/H/�Z/l/~/�//�/�$�UALRM_MS�G ?����� �/���/�/)??M? @?q?d?v?�?�?�?�?��?�?O�%SEV � �-EF�"E�CFG H�����  ��@��  AuA   Bȁ�
 O���� �O�O�O�O�O__&_�8_J_\_jWQAGRPw 2I[K 0���	 �O�_� I_�BBL_NOTE� J[JT���l�������g@�RDEFPRO�� %�+ (%�COLOCA_M�ESA_IRVI/SION�_%OVo Aozoeo�o�o�o�o�o��o�o@�[FK�EYDATA 1yK�ɞPp jG���_�������z,(����(�POINT  ]x'�)�v@NCELS��~��NDIREC�T��� EXT �STEP��*�TOUCHUǏ���ORE INFO ��C�U�<�y�`��� ����ӟ����	��-���Q�c� ���/frh/gui�/whiteho?me.pngd������Ưدꯀ{�point���0�B��T�f���  FRH�/FCGTP/wzcancel������˿ݿ�~�|�i?ndirec�(��:�L�^�p�{���nexϬϾ����������{�touchup��0�B�T�f�x���}{�arwrg�� ���������߁��)� ;�M�_�q����� ���������%�7�I� [�m����������� ������3EWi {������ �/ASew� �r������/ !/(E/W/i/{/�/�/ ./�/�/�/�/??�/ /?S?e?w?�?�?�?<? �?�?�?OO+O�?OO aOsO�O�O�O8O�O�O �O__'_9_�O]_o_ �_�_�_�_F_�_�_�_ o#o5o�_Goko}o�o �o�o�oTo�o�o 1C�ogy��� �P��	��-�?� Q��u���������ϏZj�܋�u�܏��(�s��Q�c�r�,�I���A�OINT � ]���� OOK� Tß�}�NDI�RECܟ�  CHOICE�����UCHUPG�H�s� ��~�����߯�د� ��9�K�2�o�V��������ɿ��whitehome��� ��2�D�VυĔ�poin�ߍϟϱ�����d�?i/look}���(�:�L�^�i�indirec|Ϙߪ�������g�choic���� �2�D�V�h��k�touchup��ߠ��������g�arwrg��"�4�F� X�j�a����������� ��w�0BTf x������ �,>Pbt ������/� (/:/L/^/p/�//�/ �/�/�/�/ ?׿�/6? H?Z?l?~?�?�/�?�? �?�?�?O�?2ODOVO hOzO�O�O-O�O�O�O �O
__�O@_R_d_v_ �_�_)_�_�_�_�_o o*o�_No`oro�o�o �o7o�o�o�o& �oJ\n���� E����"�4�� X�j�|�������A�֏ �����0�B�яf� x���������O�������,�>�<L�}�����u�@����q���ͯ��,�� ����"�	�F�X�?�|� c�������ֿ����� �0��T�f�Mϊ�q� �ϕ����������,� >�?b�t߆ߘߪ߼� ˟������(�:�L� ��p�������Y� �� ��$�6�H���l� ~�����������g���  2DV��z� ����c�
 .@Rd���� ���q//*/</ N/`/��/�/�/�/�/ �/�//?&?8?J?\? n?�/�?�?�?�?�?�? {?O"O4OFOXOjO|O SߠO�O�O�O�O�OO _0_B_T_f_x_�__ �_�_�_�_�_o�_,o >oPoboto�oo�o�o �o�o�o�o:L ^p��#��� � ���6�H�Z�l� ~�����1�Ə؏��� � ���D�V�h�z��� ��-�ԟ���
�� .���R�d�v������� ;�Я�����*��� N�`�r����������@�����@������	��+�=��,)�n�!ߒ�y϶� �ϯ������"�	�F� -�j�|�cߠ߇����� ��������B�T�;� x�_���O������ ��,�;�P�b�t��� ������K����� (:��^p��� �G�� $6 H�l~���� U��/ /2/D/� h/z/�/�/�/�/�/c/ �/
??.?@?R?�/v? �?�?�?�?�?_?�?O O*O<ONO`O�?�O�O �O�O�O�OmO__&_ 8_J_\_�O�_�_�_�_ �_�_�_��o"o4oFo Xojoq_�o�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t��� �����Ώ������ (�:�L�^�p������ ��ʟܟ� ����6� H�Z�l�~������Ư د������2�D�V� h�z�����-�¿Կ� ��
�ϫ�@�R�d�v� �Ϛ�)Ͼ��������h�*�`,��`���U�g�y�Qߛ߭߇�,���ߑ� ���&�8��\�C�� ��y���������� ��4�F�-�j�Q���u� �����������_ BTfx����� ���,�P bt���9�� �//(/�L/^/p/ �/�/�/�/G/�/�/ ? ?$?6?�/Z?l?~?�? �?�?C?�?�?�?O O 2ODO�?hOzO�O�O�O �OQO�O�O
__._@_ �Od_v_�_�_�_�_�_ __�_oo*o<oNo�_ ro�o�o�o�o�o[o�o &8J\3� ������o�� "�4�F�X�j������ ��ď֏�w���0� B�T�f����������� ҟ������,�>�P� b�t��������ί� 򯁯�(�:�L�^�p� �������ʿܿ� � ��$�6�H�Z�l�~�� �ϴ���������ߝ� 2�D�V�h�zߌ�߰� ��������
��.�@�@R�d�v���qp����qp����������������, 	N�r�Y������� ��������&J \C�g���� ���"4X? |�m����� /�0/B/T/f/x/�/ �/+/�/�/�/�/?? �/>?P?b?t?�?�?'? �?�?�?�?OO(O�? LO^OpO�O�O�O5O�O �O�O __$_�OH_Z_ l_~_�_�_�_C_�_�_ �_o o2o�_Vohozo �o�o�o?o�o�o�o
 .@�odv�� ��M����*� <��`�r��������� ̏�����&�8�J� Q�n���������ȟڟ i����"�4�F�X�� |�������į֯e��� ��0�B�T�f����� ������ҿ�s��� ,�>�P�b��ϘϪ� �������ρ��(�:� L�^�p��ϔߦ߸��� ����}��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� 	�������������
�������5GY1{�g,y�q�� �<#`rY �}�����/ &//J/1/n/U/�/�/ �/�/�/�/�/ݏ"?4? F?X?j?|?���?�?�? �?�?�?O�?0OBOTO fOxO�OO�O�O�O�O �O_�O,_>_P_b_t_ �_�_'_�_�_�_�_o o�_:oLo^opo�o�o #o�o�o�o�o $ �oHZl~��1 ����� ��D� V�h�z�������?�ԏ ���
��.���R�d� v�������;�П��� ��*�<�?`�r��� ��������ޯ��� &�8�J�ٯn������� ��ȿW�����"�4� F�տj�|ώϠϲ��� ��e�����0�B�T� ��xߊߜ߮�����a� ����,�>�P�b��� ���������o�� �(�:�L�^������ ����������}�$ 6HZl����� ���y 2D�VhzQ�|�>Q������ �����,�/./ �/R/9/v/�/o/�/�/ �/�/�/?�/*?<?#? `?G?�?�?}?�?�?�? �?OO�?8OO\OnO M��O�O�O�O�O�O� _"_4_F_X_j_|__ �_�_�_�_�_�_�_o 0oBoTofoxoo�o�o �o�o�o�o�o,> Pbt���� ����(�:�L�^� p�����#���ʏ܏�  ����6�H�Z�l�~� �����Ɵ؟����  ���D�V�h�z����� -�¯ԯ���
���� @�R�d�v��������O п�����*�1�N� `�rτϖϨϺ�I��� ����&�8���\�n� �ߒߤ߶�E������� �"�4�F���j�|�� �����S������� 0�B���f�x������� ����a���,> P��t����� ]�(:L^ �������k  //$/6/H/Z/�~/��/�/�/�/�/�/����+������?'?9=?[?m?G6,YO�?QO�?�?�?�? �?OO@ORO9OvO]O �O�O�O�O�O�O_�O *__N_5_r_�_k_�_ �_�_�_��oo&o8o Jo\ok/�o�o�o�o�o �o�o{o"4FX j�o������ w��0�B�T�f�x� �������ҏ����� �,�>�P�b�t���� ����Ο������(� :�L�^�p�������� ʯܯ� ���$�6�H� Z�l�~������ƿؿ ���ϝ�2�D�V�h� zό�ϰ��������� 
���_@�R�d�v߈� �ߡϾ��������� *��N�`�r���� 7���������&��� J�\�n���������E� ������"4��X j|���A�� �0B�fx ����O��/ /,/>/�b/t/�/�/ �/�/�/]/�/??(? :?L?�/p?�?�?�?�? �?Y?�? OO$O6OHO�ZO�$UI_IN�USER  ����{A��  [O_O_�MENHIST �1L{E � (�@3�(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1`�O__1_C_�'�O��N71�@BARR�A_ESTEIRAA�O�_�_�_�39X_��Eedit�BCO�LOCA�@SA_�IRVISION��_$o6oHoS_e_�A2 �Ao�o�o�o�o�Opo?,148,2�o�/AS�o�o,955o����\ov�q8�"�4�F�X��1)��o63|Q������Ϗ�����0�A����"�4�F�X�j�  ��������şן�x� ��1�C�U�g����� ������ӯ������ -�?�Q�c�u������ ��Ͽ�󿂿�)�;� M�_�qσ�ϧϹ��� ������%�7�I�[� m�ߑߔϵ������� ����3�E�W�i�{� ������������� ���A�S�e�w����� *����������� =Oas���8 ���'�0 ]o������ ��/#/5/�Y/k/ }/�/�/�/B/�/�/�/ ??1?C?�/g?y?�? �?�?�?P?�?�?	OO -O?O�?POuO�O�O�O �O�O^O�O__)_;_ M_8�O�_�_�_�_�_ �_�Ooo%o7oIo[o �_o�o�o�o�o�o�o zo!3EWi�o ������v� �/�A�S�e�w���� ����я������+��=�O�a�s�^[�$U�I_PANEDA�TA 1N������  �	�}  fr�h/cgtp/f�lexdev.s�tm?_widt�h=0&_hei?ght=10ԐŐ�ice=TP&_lines=3Ԑ�columns=�4Ԑfonܐ4&�_page=do�ubŐ1��\V) � rim#�L�   ��c�u���������$� ϯ�گ���;�M�4� q�X�������˿������%�\V� �� E�  bCFp]���ʟܝ2�����2/�-�ual ����_��"�4�F�X� j�ώ�u߲��߫��� �����B�)�f�M�`������3� E�  9��� ���*�<�N�`��� ���Ϩ��������� i�&8\C�� y������ 4Xj=���� ������� /S $/��H/Z/l/~/�/�/ 	/�/�/�/�/�/ ?2? ?V?=?z?a?�?�?�? �?�?�?
O}�@ORO dOvO�O�O�?�O1/�O �O__*_<_N_�Or_ Y_�_}_�_�_�_�_�_ o&ooJo1ono�ogo �oO)O�o�o�o" 4�oXj�O��� ���O��0�B� )�f�M����������� ���ݏ��>��o�o ���������Ο��3� �w(�:�L�^�p��� 韦�����ܯï �� ��6��Z�A�~���w� ����ؿ�]�o� �2� D�V�h�z�Ϳ����� ������
��.ߕ�R� 9�v�]ߚ߬ߓ��߷� �����*��N�`�G�����	�������������"�)��G���6� s�����������4��� ����K2oV ���������#�����$UI�_POSTYPE�  �� 	 /�U�QUICKMEN  ds�W�RESTORE �1O� � �*d�efault��  OUBLE��PRIM�m�editpag�e,COLOCA�_MESA_IR�VISION,1�0/t/�/�/;%menuH"98a/�/�/ �/?9'?4?F?X?j? |?!�?�??�?�? �?O"O4O�?XOjO|O �O�OCO�O�O�O�O_ �?_+_=_�Ox_�_�_ �_�_c_�_�_oo,o >o�_boto�o�o�oU_ �o�o�oMo(:L ^�����m � ��$�6��o�U� g������Ə؏��� �� �2�D�V�h���������ԟ�SCR�E�?��u1sc�u2��3�4�5�6��7�8��TAT`� ��M�USER�����k�s���3��4��5*��6��7��8��U�NDO_CFG �Pd����UPD�X����N�one���_IN_FO 1Q�<��0%��W���E� ��i���������տ ���:�L�/�pς�e���ύ)�OFFSEOT Td@��� {������	��-�Z� Q�cߐ߇ߙ��ϝ��� ���� ��)�V�M�_�@q�۹�����
����t��)�WORK U4�����A��S��ψ�UFRAM� ���&�RTO?L_ABRT��$�μ�ENB����GR�P 1V��Cz  A��� +=Oas��ĸ��U������MS�K  �<���N6��%4��%��)���_EVN������>�2W��
 }h��UEV���!td:\ev�ent_user\-�C7���}�YF��SP���spotweld�!C6����!�Z/�/:' �H/~/l/�/�/�/�/ -?�/Q?�/? ?�?D? �?h?z?�?O�?)O�? �?OqO`O�O@ORO�O vO�O_�O�O7_�O[_h_Z]W+�2X��F��8V_�_�_ �_ �_o�_,o>ooboto Oo�o�o�o�o�o�o �o:L'p�]�����$VARS_CONFI��Y�� FP{����|CCRG�\P��>�{�t�D�� BH� pk�a�Ce�� ��}�?����C,&Q=��ͩ�Am �MR2b��'�	}�	��@��%1: SC130EF2 *�����{�����X� �e5}�����A@k�;C�F� w�Q�[���|���������D�T����\�ϟ� �\� B���;�e�@�ǟ`����� S�����̯���ۯ� &�}��\�G�Y���E����ȿ�TCC�c�
��������pG�F�pgd���-�23456789017�?��ׁ$���4�v�Nm�� ��϶�BW�����i�}�?:�o=LA�څ �6�@�6�ͿZ���i�7����(��W���-� ]�X�jĈߚߕϳϹ� ��������%�7�I� r�m�ߨ�ߵ����� �����8�3�E�W�� ����}����������� ��/�A�S�e�w���MODE��t ��RSLT e�|k�%"zς��;� 1��d��`��SELEC��c�}�	IA_WO�P�f �� >W,		�����>�G�P ������RTSYNCS�E� ��$�	#WINURL ?*ـ�;\/n/�/�/��/�/�uISION�TMOU���A# ���%�gSۣ��SۥP�� �FR:\�#\D�ATA\�/ �߀ MC6LO�G?   UD�16EX@?\�'� B@ ����2T1Gabri�el_Faria�k?P5�?�?������ n6  ����GV�2\� -�|�5��   ���Z�@U058TRACINj?��*B{Rd_C�p��D #A`{2��'$�"��h#� (�kI�Mw��O �O�O�O�O1__U_C_�]_g_y_�_�_�_�(SKTA� i��@���o0oI:$obo�%_kGE�j#��~@� �
�\��btgH�OMIN�kS����`�2,,���CWǖBveJMP�ERR 2l#�
  QoI:��"� 4Fwj|����������&%S-_g0RE�m�^۴�LEXdn�1�-ehoVMPHA�SE  �e׃�BޱOFF _E�NB  �$V�P2�$oSۯR��x�c C;�@ ��@�;���?s33'D*AA��]� �P�0ޱ�`r}�XC ��܅���\A-۟E ������#� 5�������������}� ���������c�X� ��A�����ϯ�+�� ߿��M�B�q���x� �Ϲ���Ϸ������� 7�I�;�m�b�)ߣ�E� �ߡ߳�����3��� W�L�{ߍ��ߑ��� �������/�$�6�e� W���c�y��������� �����O���?M _q������� '9�=7Is� �����/m�/%/3/E/s�TD__FILTE�`s�kg �x2�`��� �/�/�/�/�/	??-? ??Q?�6�/~?�?�?�?��?�?�?�?O OoiS�HIFTMENU� 1t}<5�% 5�~O)�\O�O�O�O�O �O�O�O'_�O_6_o_�F_X_�_|_�_�_�_�	LIVE/SN�AP�Svsflsiv���_�z`/ION ҀU
`bmenu&o+o�_�oP�oV"<E�uz��4IkMO�v���zq��WAITDINEND  �ec��b��fOKوOUT��hSDyTIM.du��o|G�} #�{C�zb�z�x�RELE��ڋxT�M�{�d��c_A�CT`و��x_D?ATA wz����%  EGA_B�ARRA_EST�EIRA�o6Ex�R�DIS
`E��$�XVR�ax�n��$ZABC_GRoP 1yz���� ,�2̏.MZ�D��CSCH�`zd���aP@�h@�IP�b{'����şן�[�MPCF__G 1|'���A0�r�8��� �}'���p�s� 	|(���  <l0�  ��  ����5�>�����?��5�`���?5�U������C�Tp���1V�>w�@3�>�?|�/�Q���6 `��@Q�>���`���� ��˯ݯ����o�p��w���� /��C3����"��3��˿ݸĸ� �	��1�?�i���'�9�0?�Q��	��`�~����_CYLI�ND~!� ��� ,(  * .�?ݧ+�h�Oߌ�s� ��������(�	� x�-��&�c�߇�� ������j�P����)���~�_�q��� �2�'��� �&���� ������&��I��cA���SPH�ERE 2��� �������A� T/A��e�� ����/N` =/�a/H/Z/�/��/��/�/�ZZ� � �f