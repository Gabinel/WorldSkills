��   T�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ������DMR_SHF�ERR_T  � $OFF�SET   w	��/GRP:�� $MA���R_DONE � $OT_M�INUSJ  	�sPLzdCOU=NJ$REFj��PO{��I$�BCKLSH_S�IG�EACH�MSTj�SPC��
�MOVn ~A�DAPT_INE�RJ FRIC�COL_P,MGRAV�� �HISIDSP|k�HIFT_7 -O �Nm��MCH� S�AR�M_PARAO� dcANGo zy2�CLDE7��CALIBD~n$GEAR�=2� RING���<$]_d�RE�L3� 1  �	��CLo:o � �AX{ � $PS_�T�I���TIME� �J� _CMYD��"FB�VA >�&CL_OV�� oFRMZ�$DE�DX�$NA� =%�CURL�qW���TCK�%��FMSV>�M_LIF	���'83:c$�-9_09:_��=�%3d6W�� �"�PCCOM,��FB� M�0�oMAL_�ECI��P:!o"DTY�kR_|"�5:#�1E�ND�4��o1� l5M�P P�L� W ��S�TA:#TRQ_MH��� KNiFS� �uHYsJ� hGI�JI��JI�D��$�A{SS> ����A������@VER�SI� �G�  0��AIR�TUAL�O�AS �1�H }��� 	 �� \_G_�_k_�_�_�_�_ �_�_�_"oj�ABo0o� ��������DP� f����Wo�o+oUl�o@�o�o�o�o�k;�Ar*gyd���d�������=L̙���?����@�=�b�t����������Ώ�����(�{ �US�a�K����D  2���ğ֟���@��0�B�T���<�� ~�������Ưد����� �2�D���Pr�( �x����������� Ͽ���>�)�b�Mϰ��qϖϼ��$4 �12\���E��� F@ ��5W�ś�ߗ� @�M�Aߚ�h�z�e� ��9�K߅���߈��� �9�$�]�o��X�S�X�\�X�,���� ��������������,���%���345678901G�O�t�x�q��� m�����������D� }���z�H��lZ |�����.� �2 Vh��� �n@���/r �U/���//�/�/ �/�/8/	??n/�/N? <?r?`?�?�?�/�?"? 4?�?�?O8O&O\O�? �?�O�?�?�OFO�O�O �O"_xOI_[_�O_�_ |_�_�_�_�_>_ob_ t_�_�_Boxofo�o�_ o�o(o:o�o, <b�o���oP� ����(�~O�� �.� �������܏2� D��h�z�H�Əl�Z� |�����ɟ۟.���� ��2� �V�h������ ��n�@�¯����r� ��U������������ ���8�	��n�пN� <�r�`ϖϨ�����"� 4Ϯπ��8�&�\�n�`}��ϕ����%�B����8��$PLCL�_GRP 1S��� D�?�  ��� ;��_�J��n��� ���������%��