��   �;�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_CPC�_T 4 $�COMMENT �$ENAB�LE  $M�ODJGRP_N�UMKL\  $UFRM\~] _VTX M ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�? �ELAY_T�IMJSPEED�_CTRLKOV�R_LIM? p JD� L��0�UTOO(i��O��&}S. � 8J\TC�u
!����\� �jY0  � ��CHG_SIZ��$AP!�E.�DIS�]$!B�C_+{#s%O#J�
p 	]$Jd#� �&s"��"{#�)�$�'�_S}EEXPAN#�N�iGSTAT�/ DFP_�BASE 5$0K$4!� .6K_V7>H73hJ- � }�\7AXS\UP�LW�7���
0c5r �< w?�?�?���?�?�//	7E�LEM/ T 1�&B.2NO�G]@�%CNHA�DF#� _$DATA)he0  PJ�@� 2 
&PN5 �� 1U*.n   _VSiSZHbRj0jR(�VyT(��R%S{TROBOT��X�SARo�U�V$CUR_��Rj�SETU4"	 ��bAISP_MGN��INP_ASS e#�PB!� `CiH�7�7`e�.fXc1�C�ONFIG_CH�K`E_PO* }dS/HRST�gM^#/e�OTHERRBTF�j_G]�R�dTv ��ku�c)&T1r
�0R HLH�d� 0  �lt<Ne'AVRF!YhH^t�5�1� �r�W�_A$Rdv�TPH/ (@G%Q�Q�Q3wwBOX/ 8�@ F!�F!�G �r{�z�TUIRi@ c ,�F�pER%@�2 $�p [L�_SF�!�ZN/  IF1(@�p��Z_�0��_�0wu0  @��Q7yv	
��~ ��$$CL`  O������Q���Q��VERSIO�N��  �0��IRTU�AL���' 2 ��Q  (�p���&@>�m��P��������������Ғd��Cz  0����A��� l���������Ɵۯ� ��� �2�D�F�h�}� ����ԯſ�����
� �.�@�R�d�fϋϚ� ����п���ώ��*� <�N�	�rχߖϨ�b� �Ͼ�����&�8�^� \�n߃��߶����� ����"�4�F�X�m� |������������ �0�B�h�Vx�� ���������� ,>Pbw��� ����//(: L�`/��/��� �/�??$/6/H/Z/ l/�?�/�?�/�/�?�/ �?O#O2?D?V?h?jO �?�O�?�?�?�O�O_ _.O@OROdOvO�O�_ �_�O�O�_�O	oo�_ <_N_`_r_-o�_�o�_ �_�o�_�o)8oJo \o�o�o�o�2�o�o ��o�%�4FXj |���������� ��!�3�B�T�f���z� ������ҏ����� /�>�P�b�t������� ��Ο������+�=� L�^�p��������ʯ ܯ���'�9�H�Z� l�~����ϴ���ؿ� ���#�5�G�V�h�z� �ώ߰��������� ��1�C�R�d�v߈ߚ� �߮�������	��-� ?���`�r���Q��� ��������;M \�n����������V ����"7IXj |������� �/E/W/fx� ��/��/��/? ,/A?S?b/t/�/�/�/ �?�/�?�/?O(?=O OOaOp?�?�?:O�O�? �O�? OO'_6OK_]_ lO~O�O�O�O�_�O�_ �O_#o2_GoYokoz_ �_�_�_�o�_�o�_
o @o1 Ugvo�o�o �o�o�o��-� <Q�c������ u�����Ώ8�*� _�q�������ʏȏڋ��$DCSS_C?SC 2����Q  AP����:�܉d
� k�.���R���v�ׯ�� ��Я1���U��y� <���`���ӿ������ �޿?��c�u�8ϙ� \Ͻπ��Ϥ������ ;���_�"߃�Fߧ�j� ���ߠ����%���I� �m�0���f���������GRP 2��� ����	 ҟS�>�w�b������� ��������=( aL�p���� �� K6o Z�~����� �/5/ /Y/D/}/h/ �/�/�/�/�/�/?�/ 
?C?.?g?R?�?�?�? z?�?�?�?�?O-OO QO<OuO�O�OdO�O�O �O�O_�O_;_&___ q_�_N_�_�_�_�_�_��_�_%ooIo��_GSTAT 2��~%��< ���F��>�:Z��L?!h�>��l�3�����¿M���5?>���Ġ^�A;}���8`<�e8�(�����4��Z.O#^�?�`�a��`~�a<�g�������ft_�����?_&׸���]q>p�i=W�����D��� z�]��1R��?8��a8�����-��/�PrMp=��d����D&��� y:��-hp߿8�����zdu�?�뺅�h�:���>��Ė[7B�!>~x{ї?53�`�ٿ�p:��غ����8�v?M��pB��o�o �o y��<�N���0�z� ��f���Љ�i�a-i ��+k y �.��&�H� v�\�~��������ȟ ڟ��*���Z�l���x� ��|���د���.�� B��J�0�B�d���x� ��ȿ���������� F�H��Ϻ�tϾ���������͵����?�6<�R���a5��t��j߷��P4�޿��5@�K�C�"D)���m�<rE�?���5a����1�~ɯ�apѼm��a@���C��,ͼ�Mq�YR?���� gʿ�ٿYe������ó`�C�� y��Q�>��� ?r��;�q�<rDN�����eњ��r�p������Ǹ����Cw�ް�ڌ�-��}���:�e�� ��p��pK&����@�MCĿڑDB�� y<�p]�?�)<��MJ���<pK�9��/5��}�I�0�O�F�(�:� L����������� ��� �V�h��Pϒ�dϪ� ����������F ,^|bt��j� �8��<N(r �z������� ��,//4/b/H/Z/ |/�/�/�/�/�/�"? T?X?j?D?�?�?z? ���P�b�t߆ߘߪ� ����������(�:� L�^�p��O�?�?�?�? t_�_|?�_�_�_�_�_ o��/.o ?FodoJo \o~o�o�o�o�o�o�o �o2`?�� �_����� �o dJ�xB�d���x��� ȏ��Џ������F� ,�N�|�b�(������ �����*�<��4_F_ �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O _~�`�r�����"� �.�X�2�DώϠ�:� ���Ϝ��� ������ H�.�P�~�dߖߴߚ� �����ߢ�,�>�p�*� t��`���� ��� ��� �.��6�d�J� l��������������� ����Z��F�� |���п⿈��� ����Я�����*� <�N�`�r�������/ � ��/�/��/ �/�/�/*?<?��$f? 8~?�?�?�?�?�?�? �?O O2OPO6OHOjO �O>�O�O?�O_"_ �OF_X_N?�O�_�Oz_ �_�_�_�_ o�_o6o o.oPo~odo�o�o�o `_�o(_�o,>b tNl/~/$6HZ l~������ �/ /2/D/���� �VH�Z�Pf���j� |�Ɵ؟r_�o��o� 8��0�R���f����� ��ί�ү��4��o d�v���b�������� ���8��L��8�f� L�nϜςϤ��ϸ��� ��� �"�P�6����� Ŀ~����ߴ������ �������� ,�>�P�b�t������� ��Ώ��R�4�F�X��� ������,b t�\ߞp߶�� ��$R8j �n���v� // D�H/Z/4/~/�/� ��/��/�/?�/
? 8??@?n?T?f?�?�? �?�?�?�?�/.O`/O dOvOPO�O�O�O���� \�n��������� �����"�4�F�X�j� |��_�O�O�O�O�o�o �O�o�o�o�o�o�/ �?:ORpVh� ������$�
� �>�l�O�����o�� ���Џ�,�"p�V� ��N�p�������ԟ�� ܟ
���$�R�8�Z� ��n�4�ʯ���� ����6�H�V��$DC�SS_JPC 2�@�Q �( DMP���� ����P��ۿ����� ���Y�(�g�Lϡ� p��ϔ��ϸ����1�  ��g�6�H�Z߯�~� �ߢ��������?��  �u�D�V�h����� �����)���M��.� p���d�v��������� ��7[*N �r�����! �/i8�\� ������//� /"/w/F/�/j/�/�/ �/�/?�/�/=??? 0?�?T?�?x?�?�?�? �?O�?�?8O]O,O>O �ObOtO�O�O�O�O�O #_�OG__k_:_L_�_ p_�_�_�_�_�_��h�Sq�u�L�_Uooyo��dDo�oho�o�o �o�o�o1�oU y@Rd���� ���?��c�*��� N���r�����󏺏̏ ޏ��M��q�8���\� ����ݟ���ȟ%�� ���Y��F���j�ǯ ��믲��֯3���W� �e�B���f�x����� ������A��e�,� ��Pϭ�t��ϘϪϼ� �+���O��s�:ߗ� ^߻߂��ߦ����� ��K��$�6�H��l� ���������5��� Y� �}�D�V�h����� ��������C
g .�R�v��� ����Qu< �`����/��&dMODEL 2�3kx��
� <�c (  �z(�/g/y/ �/�/�/�/�/�/�/D? ?-?z?Q?c?u?�?�? �?�?�?�?.OOO)O ;OMO_O�_�OY/�O�O _�O�O<__%_7_�_ [_m_�_�_�_�_�_�_ �_8oo!onoEoWo�o {o�o�o�o�o�o�O�O �O�o|�oew� �����0��� +�=�O�a�������� ��͏ߏ���b�9� K���3Es����m� ۟����#�p�G�Y� ��}�������ůׯ$� ���Z�1�C�U�g�y� ��ؿ����ϩ���� ��h��Q�cϰχϙ� �Ͻ��������d� ;�Mߚ�q߃��ߧ߹� ������N�%�7�� �1�C�q��Y����� &����\�3�E�W�i� {������������� /A�ew� ��������� �=O�s��� ����/P/'/9/ �/]/o/�/�/�/�/? �/�/:??#?5?�? /]?o?�?�?�?O�? �?HOO1OCO�OgOyO �O�O�O�O�O�O�OD_ _-_z_Q_c_�_�_�_ �_�?
o�?�_�_Ro)o ;o�o_oqo�o�o�o�o �o�o<%7I [m������ ���!��_��oI� [�ȏ������Տ��� ��/�|�S�e����� ������џ�0��� f�=�O�a�s�����m� ������ѯ>��'�t� K�]�o��������ɿ ۿ(����#�p�G�Y� ��}Ϗ��ϳ�����$� �������5�Gߴ� /ߝ߯�������2�	� �h�?�Q�c�u��� ����������)� ;�M���q�����k�}� ����*��%7I [������ ��\3E�i {����/�� F/����!/3/�//�/ �/�/�/�/?�/?T? +?=?O?�?s?�?�?�? �?O�?�?OPO'O9O �O]OoO�OW/i/{/�O �O�O�O_^_5_G_�_ k_}_�_�_�_�_o�_ �_Hoo1oCoUogoyo �o�o�o�o�o�o�o�O V�O1u�� ��
�����)� ;���_�q��������� ˏݏ�<��%�r�I��[�m����$DCS�S_PSTAT ����ӑ�Q    ��� � (��+��O���t� r�Ԑ�������������ӕ௎�կ��ĔSETUP �	әBȖ��� ��8�R�ͬs�b����������T1SC 2i
+�����Cz�������صCP R-�D�DLj� |�>�ϲ��ϓ����� ���0�B�T�#�xߊ� Yߛ����ߡ����� ��>�P�b�1���� y��������(��� L�^�p�?��������� ��������$6Z l~��Vϫ�D� ��);Mq ��d����/ /�7/I/[/*//�/ �/r/�/�/�/�/?!? �/?W?i?8?�?�?�? �?�?�?�?�?O/OAO OeOwOFO�O�O�O� �O�O_�O+_=_O__ s_�_�_f_�_�_�_�_ oo�_9oKo]o,o�o �o�oto�o�o�o�o #�oGYk:�� �������1�  ��g�y�H������� �����	��O-�?�Q� ؏u�����h���ϟ�� ����;�M�_�.� ������v�˯ݯ���� �%���I�[�m�<��� ������ٿ���̿!� 3��W�i�{�Jϟϱ� �ϒ��������/�A� S�"�w߉��j߿��� ��������=�O�a� 0����x������ ��'���K�]�o�>� ���������������� #5Yk}L� ������1 Cgy�Z߯� �Z�	//�?/Q/ c/2/�/�/h/z/�/�/ �/??)?�/M?_?q? @?�?�?�?�?�?�?�? O%O7OO[OmOONO �O�O�O�O�O�O�O�O 3_E__i_{_�_\_�_ �_�_��_oo�_Ao Soeo4o�o�ojo�o�o �o�o+�oOa sB��x��� ��'�9��]�o��� P�����ɏ�����Ώ #�5�G��k�}���^� ��şן�������_ C�U�ܟ6�����l��� ӯ寴�	��-���Q� c�u�D�����z�Ͽ� �¿�)�;�
�_�q� ��RϧϹψϚ���� ��%�7�I��m�ߑ� `ߵ����ߨ�������3�E�W�&��$DC�SS_TCPMA�P  ������Q @� .�.�.�T.���.�.�.�U.�	.�
.�.�U.�.�.�/�W  .�.�.�U.�.�.�.�.�.�.�.��.�.�.�.� �.�!.�".�#.�$�.�%.�&.�'.�(�.�).�*.�+.�,�.�-.�..�/.�0�.�1.�2.�3.�4�.�5.�6.�7.�8�.�9.�:.�;.�<�.�=.�>.�?.�@�u�UIRO 2.��������� ������,>P bt�������-���-��Q cu������ �//)/;/M/_/q/ �/�/2�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O�/ 3O�/WOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_&O�_q�UIZN 2��	 ����� oo $o*��_Rodovo9o�o �o�o�o�o�o�o* <Nr��Y� �����&�8�� \�n�=�������ȏ�� ����ߏ4�F�X�� |�����o�ğ֟蟫� ��0���T�f�x�;� M������������_~x�UFRM R�����81�^�p� /����ʿܿ�� � ��6�H�#�l�~�Y� �ϴϏ��������� � 2�I�V�h�ߌߞ�y� ���߯���
���.�@� �d�v�Q����� �������*�A�N�`� �����q��������� ��8J%n� [������ "9�FX�|�i �����/�0/ B//f/x/S/�/�/�/ �/�/�/??1(?P? b?=?�?�?s?�?�?�? �?O�?(O:OO^OpO KO�O�O�O�O�O�O _ _)?;?H_Z_�O~_�_ k_�_�_�_�_�_�_ o 2ooVohoCo�o�oyo �o�o�o�o
3_@ R�ov�c��� ����*��;�`� r�M�������̏ޏ�� ��+8�J��n��� [�������ǟ���ٟ "�4��X�j�E����� {�į֯������