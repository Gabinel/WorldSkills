��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ��!PCOUPLE�,   $�!PPV1CES C G�1�!�� A> �1	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q�RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Nb_OPT�2 �� ELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1� UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t���MO� �sE 	� [M�s��2�wREV�BILF��1XI� %�R 7 � OD}`j��$NO`M��!b�x�/��"u�� ����4AX��@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC���a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���OR4@BIGALwLOW� (KtD2�2�@VAR5�d!�A}#BL[@S �� ,KJqM�H`S�pZ@M_O]z����CFd XF�0GR@��M��NFLI���;@U�IRE�84�"� SgWIT=$/0_No`�S�"CFd0M�� �#PEED���!�%`���p3`J3tV�&$E�..p�`L��ELBOF � �m��m�p/0��CP�� F�B�����1��r@1J1E_y_T>!Բ�`���g���G� �>0WARNMxp�dp�%`�V`NST� �COR-rFL{TR�TRAT �T�`� $ACC�qM�� R�r$OcRI�.&ӧRT�sSFg�0CHGV0I�p�T��PA�I{�T�!��� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8��9/C���x@�2w @� TRQ���$%f��ր����_�U������Oc <� ����Ȩ3�2^��LLECM�-�MULTIV4�"$���A
2q�CHILDh>�
1��Oz@T_1b�  4� STAY2�b4�=@�)2�4����@�� | 9$��T�A�I`�LE��eTO���E��EXT���ᗑ�B�᎞22�0>���@��1b.'��B 9�A�K�  �"K� /%�a��R���?s��?�O�!M��;A�֗�M8�� 	�  =�I�" L�0[�� �R�pA��$JOB`B���������IGI�# dӀ����R� -'r��A�ҧ_��`�n�b$ tӀFL6��BNG�A��TBA � ϑ�!��
/1�À �0���R0�P/p ,����%�|���Bq@W�
2JW�_RH�CZJZ�_zJ?�D/5C�	�ӧ���@��;�Rd&A������ȯ�qGӨ�g@NHANC��$LG/��a2qӐ� ـ�@��A�p� ���aR���>$x��?#DB��?#RA�c?#AZ�t@�(.�����`FCT����_F࠳`�SM��!I�+lA�% ` �` ���$/�/�@���[�a��M�0�\��`��أHK��A�Es@͐�!�"W��Nz� SbXYZW�`$�"����6	�������'  . I�I��2�(p�STD�_C�t�1QA��U+STڒU�)#�0U�[�%?IO1���� _Up�q�* 1\��=�#AORzs8B�p;�]��`O6  RSY�G�0�q^EUp� H`G�� ��]�@P_XWORK�+^�?$SKP_�p��DB�TR�p , �=�`����Z �m�OD3��a _C`"�;b�C� �GPL:c�a�tőS�D�W�3Bb����P�.�&�DB�!�-�B A{PR��
�DJa3��. /�u���.����LuY/�_�����0�_�� ��PC�1�_���r~�EG�]� 2�_���I�
!.��R3H� $C��.$L8c/$uSނz IkgINE�WA_D1%�ROyp�������`�q�c7 t@�fPA��~�RETURN�b.��MMR"U��I�;CRg`EWM@�/SIGNZ�A ����e� 0$P�'�1$P� m�	2p�p'tm�+pD�@ �'�bdNa)r�GO_AW ��h@ؑB1@CSd��(�CYI�4���`1Pw�qu��t2�z2�v�N�}��E}sDE�VIs` 5 P7 $��RB���I�wPk��I_B�Y���"�T7Q�tH�NDG�Q6 H�4��1�w��$DSBLC��o��vg@��4sPqL��7O�f@�]���FB���FE�ra8�ׂ�t}s���8�> i�T1?���MC�S���fD �ւ[2H� W��EE���%F���Ů@q����9 Tx�p��x�NK_N:�Ԅ���U��L�wHA�vZ��~�2���P�~r�q7: �=MDLn���9�ጂٱ h����!e����J��~�+����,�N�D����3��ՒG!a�qSLAd�7;  ��INP��"������}q_ �4<�0�6`C� NU�� � D�Lק� h�_ S)H!�7=M��q⑄��ܢӢ��������>P +$ ٰ�٢��^��^�Y�FI B\��Ă���'A	'AWl�N�TV��]�V~�X�SKI�#T���a�ۺ$�T1J�3:3_�P��SAFN���_S}V�EXCLU��*N@�DV@L��@��Y����S�HI_V�
0\2PPLYPR�o�HIM�T�n�_M�LX��pVRFY�_�Cl�M��IOC�UC_� ����O�q�LS�0v�FT%4Q�����@�P�E$�t��A��CNFt�6եu��pm�4ACHD�o����6��AFC CPlV��TQ����_�� ?`�@TA�@�0L@� )�8��N���]� @����T��T! S����te@{R�A DO�� w23���!n��	_1�#�H!�f��΀�K��B�2��MAR�GI�$����A �̔_SGNE�C;
$�`�a^aR0 ��3��  B��B��ANNUN�P?����uCN@�`%0��`��� ����EFc@]I�RD @Q�F���4OT�`�sFT�`HR,Q��CQ�pEM��NI|RE�����AW���DAY=CL�OAD�t;T|�<S5�}�EFF_AXIJ��F`1QO3O��|�S�@_RTRQE�eG����0RQj��Evp ���F��0f�R0 �te��AMP�E<� H 0�`œ^�`LDs�DU�`���B;CAr� I?�`�N ErIDLE_�PWRI\V!n0V��wV_[ ꐅ �D�IAG�5J� �1$V�`SE�3T Ql�e��Pl�f^E_��j�VE� �0SWH�q(�� C2�Gn�O�HxPPHk�I	RAl�B�@�[��a �bk��w3�O � ��v��I�0 �p�RQDW�MS�-�%AX{6j�LIFE�@�&�MQy��NH!Q%��F#CD����CB0�mpN$�9Y @D1FLAl���3OV0]&HE��l��SUPPO�@u��y��@_�$��!_XP83�$gq�'Z�*W�*�B1�'T�#`�k2XZ�áj�Y2D8CY`T@�`N����f�� �C�k�̒ICT�A�K `�pCACH�ӫ�3����I�z�bNӰUFFI� \��@��;T��<S�6OS�@MSW�5L� 8	�KEYIMAG�cTMLa��*A�x�&E���B��OCVsIER-aM ���BGL����y�?�G 	U�@�П4N�m:�ST�!�B P�D,P�D��D��@EMAI䐔a��sP^s�FAUL|RObB�c�� spUʰ�`X �DT'`E�P< �$S�S[ � ITw�BUF�7y��7r�tN[�LSUB1T��Cx�o�R�tRSAV|U>R'c2�\�WT���P�T�*`S�n�_1PbU���YOT(�bK��P��M��d����WAX��2��XX1P��S_GH#
�p�YN_���Q <���D��0���M��� T�F�`�|�\�DI��EDT�_Pɰ:�R��b�GRQM�&��Jq�a�1׀���Fs� S (�SVqpB��4�_����a��T� ��@���B�SC_R]1IKU'r��$t���R"A#u�H�aDSPd:FrP�lyIM|S as�qz��a� U>w� 4<1%sM�@IP��s��0`tTHb0ЃTr2��T`asHS�cCsGBSCʴq0� V������S�_D��CONVE�G���b0$^v1PFHy�dCs�`�&aVSC���sM�ERg��aFBCM�Pg��`ET[� mUBFU� DU%Pb�D�:12�CDWy�p�P�C�`R��6�:�AV� ��� ���P�ъ�C����w��Q��`��WH *�LƠ�Cc�W��� �Y�賂��р�q�@|���A��7}��8}�9}�H ���1���1��1��1��1�ʚ1ך1�1�2R��2����2��2��U2��2ʚ2ך2�U2�3��3��3�����3��3��3ʚ3*ך3�3�4��Ka'EXT[�X[b�H�``t&``z�k`˷$��� �FDR�YTPV��RK"�	��K"REM*F���]"OVM:s/�A�8�TROV8�DTl�PX�MXg�IN8�8� W��INDv�["!
�ȕ`K ^`G1a��a��@Q%7Da�R�IV��u"]"GEA-R:qIO.K(�[$N�`���,(�F@� >\#Z_MCM<0K!��F� UT���Z� ,�TQ? �b�y@t�G?t�E |ј>Q�����[@�Pa� R�I�E��>SETUP?2_ \ �@=S#TD	p<TT����p����q>RBACUbG] T��>R�d)�j�%C�E��0��IFI���0��i�{�4�PT�T�AFLUI�D�^ Ђ gHPUR �gQ�"�r�a�4P�+ I�$��Sd�k?x��J�`CO�P��SVRT��N�x$�SHO* ��CAS�S��Qw%�pٴBG_%��3���<�FORC�BZ�^o�DATA��_�BKFU_�1�bb�2�a�ge,m�b0��` �|��NAV	`)������$�S�Bu#?$VISI���2SC	dSE������V��O�$&�B�K�� ��$PO���I��FM�R2��a  ��	��`#��@&�8�O� (�_��9��+IT_^�ۄ�)M�����DGC{LF�DGDY�LD����5Y&��Q$RY�M됇CbN@{	? T�FS�P�D�c P��W�cK �$EX_WnW1P%`]��"X3�5�s�G+�d ���ָ�SWeUO�DE�BUG��-�GRt��;@U�BKU���O1R� _ P�O_ )�����M���LOOc>!SM E�Rq��u _E e � ���@�TERM`%fi'O�ORI�ae gi%�y�SM_�`>Re h�i%V�(ii%3U}P\Bj� -��F�e��w#� f��yG�*ELTO�A9�bF�FIG�2�a�_���Ў$�$g$U;FR�b$�1�R0օ� OT_7F�TqA�p q3NST�`�PAT�q�0�2PT�HJ�ԀE�@�c3ART�P'5�Q��B�aREL�:�aS�HFT�r�a�1�8_���R��у�& � $�'@i�
����s@b�SHI�0�Uy� �QAYLO�p�Oa�q�����1����pERV��XA��H��m7��`�2%�P�E3�P�RyC���ASYM�a���aWJ07����E �ӷ1�I��ׁUT�` Oa�5�F�5P�su@�J�7FOR�`M  �O!k]��5&0�0L0���HOL ;�l �s2T����O�C1!E�$�OP��qn���H$�����$��PR^�f�aOU��3e���R�5e�X�1 �e$7PWR��IMe�BR_�S�4�� �3�aCUD��p�Q�dm���$H�e!�`AD+DR˶HR!G�2�a��a�a���R��[�n H��S����%��e`3��e���e��SEl�� HS�MNu�o���Pªq��0OL�s߰`ڵ�I ACRO��&1��ND_C�s��Afd�K�ROUP��R_�В� �Q1|�=�s ���y%��y-��x���y���y>�=A��Ҁ��AVED�w-��u,<&sp $���P�_D�� ��'rPR�M_��HTT�P_�H[�q (�ÀOBJ��b �$˶LE~3�P��\�r � ���ྰ%_��TE#ԂS�PIC��KRLPiHITGCOU�!��L�� �PԂ������PR��P�SSB�{�JQUE?RY_FLAvs�@_WEBSOC��G�HW�#1��s�`}<PINCPUPr��O���g�����d�t��O��IO�LN�t 8��R���$SL!$INPUT_U!�$`��P M ֐SL.���uᐁ��2�.��C��BL�OG֐a�F_AS=v�$a�ʷy�NA��bb41�����Z@HYʷ�����#qe�UOP:w `v�ϡ˶�¡�������"`PIC`����� �	�H�IP_ME���v�x Xv�IP�`PrR�_N�p�d����Rʳp��QrSaP �z�C��BGPq� ��M�Av�y lL�@CTApB��AL TI�3UfP_ ۵�0�PSڶBU_ ID � 
�L � `�; ��L��0z)�����ϴ�NN�_ O��I�RCA_CNf� �{ �Ɖ-�CYpEA������� �IC�ǫ�tpR�=Q�DAY_
��NTVA�����!��5�����SCAj@��CL��
����
���v�|`5�VĬ2b�l�N_�PACV�n�
���w�})� T��S�����
��e����T� 2| c��� �v�~��֣�ذLAB1��_ �חUNIX��ӑ I�TY裪��e���p�� ��<)���R�_URL���$A;qEN ���s`vs�TeqT_U���iJ��X�M�$���E�ᒐR祪�� A��,���JH���FL�y��= 
���
�wUJR|U� ���AF�6G��K7��D>��$J7�s��J8B*�7���3�E�7���&�8\�)�APHI�Q4�y�DkJ�7J8R��L_K�E'�  �K�͐LMX� � �<U�XRi�����WATCH_VAZqxu@AំFIEL`�b�cyn���:� � bu1VbwPCTX�j�Y �LGE�߄� !��LG_SIZ΄�[8XZm�ZFDeIY p1!gXb ZW �S `�8�m��� ��b ��A�0_i0_�CMc3#�*'F Q1KW d(V(Bbpo pm�p� |Io�1 p�b pW RS��0 7 (n�LN�R��۠�DE6E�3����c�i���PL�#�DAU"%EA`q�͐�T8". GH�R�:�a�BOO�a��� C��F�IT0V�l$A0��RE���(GSCRX����D&�|ǒ�qMARGI4� Sp�,����T�"�y�	S��x�W�$y�$���JGM7MNCHLt�y�FN��6K@7�r�>9UFL87@L8F�WDL8HL�9STPL:VL8"�L8s L8�RS�9HOPh;��C�9D�3R��}P�'IU h�`4�'�5$ ��S2G09�pPOWG�:�%`�3,64��N9EX��TUI>5I� �ӌ������C3�C<0'�@,�o:��&�@�!Naq�vcANAy��Q�A�I]�gt7Ӝ�DCS����cRS�cRROXXO"dWS�ÂRoXS{X�(IGNp 
Ђ=10 ܰ�[TDEV�7LL ��Ԑy��C �	 8�Tr$f/蛒�Ĵ��3A�a�	 �W�萦�Oqs�S1
Je2Je3Ja��BSP�C � �ƋG`-T ��%��Q�T�r@�&�E�fST�R9 Y�Br�a �$E�fC�k�g��f	vB��DB� L�����  ��u�xs뀔�g�q�jt�jd�$_ � �[��w�#Ӡ �s �{MC�� ����CLDP᠜�TR�QLI ���y�tFAL���rQ��s5�D���w~�LD�u�t�uO�RG���1�RESERV��M���M��Œ��s��� �� 	�u�5�t�uSVH��p��	1�����RCLMC��M�_��ωА��: MDBG�h�I����$DE?BUGMAS�������U�$T8P��E�F�d���MFR�QҤ� � ~K	HRS_RU4��bq��A��$EFR3EQ6u!$0YOVER�k��f��PU1EFI�!%Gq�� �aY�z�ǐ \����E�$9U�`��?��
�SPSI`��	��CA ���ʲ�σUY�%��?( 	��MIS�C�� d��aR5Q��	��TB� �c ���A��AX����𑧪�EXCESHg�!qd�M�H�9��u���`@c�S}C�` � H����_����������
b�KE��+�� &�{B_, FLICBt}B� QUIRE C�MOt�O��얩qL:dpMD� �p{!���5b���r�ND!��I����L ��D;
$INAUT�!
$RSM�ȧPaN�b�C�$L��PSTLH� 4nU�LOC�fRI"�v�eEX��ANG.R�.�W�ODA]��bq��� ���MF0 ����icrO@mu����$�SUPvv��FX��IGG! � �O�cs��#cs
F ct��ޒ�b5��`E��`�T�5�tC��g�TI���7b�� M����� tZ�MD���) ��XP��ԁ��H��.���DIAa��Ӻ�W��!��0af���D@#)��O�㥀��� �CUp V	���.��֡O�!_��� ��{`�c������� |�P|��0� ��P�{�KEB��e-$qB��o�=pND2ւ�����2_TXltXGTRAXS������LO: ���������C�.�&��[�RR2h���� -�!A�� ?d$CALI����GFQj�2F`RIN�bn�<$Rx�SWq0ۄ���ABC�ȇD_J��{�q��_�J3��
��1SPH, �q�P����3��(H�9pq�#J�34n���O�QIM�M�CSKP�zb7?SbJ+�M�Qb�y8����_AZ��/��EL�Q.ցOC�MP��N�� RTE�� �1�0 ����1��@ ZScMG�0����JG�p�SCLʠ��SPH�_�PM��f��q��u�RTER��n��Pk�_EP�q�`A0� �cM��DI�Q�23UdDF  쀐�LW�VEL��qINxr�@�_BALXP.��Y/�J���'$���IN���]�C�9%�".��8!6p_T� �@F%a"�j`^$��k)��"pDHʠ��\�9`$Vw��_�A�$=��~�&A$�����R6�]�H �$BEL� |m��_ACCE�� 	8�0IRCi_�q�@�NT���c$PSʠ�rL���M4�s9 .7���GP/6��9�7$3�73S2T�͡_Ga�"�0�1���8�1_MG}�D1D�1�~�FW�p��`3�5$32�8DEK�PPABN[7ROgEE�2KaBO�p��Ka��1�$U�SE_v�SP��C�TRTY4@� �� <qYNg�A�@�FR ��ѢAM:�N�=R�0O8�v1�DINC(���B�4���GY��ENC�L��.�K12��H0IN�bIS28U���ONT�%NT2c3_�~�fSLO�~�|P��Iذ��V�@�$��hpU#�CQ MVMOSI�1<�[���1��M�PERCH#  �S��� �W�� �SlщR��l����EH�0�0PAS2EeL�D P7�ONUЉZ�f�VgTRK�RqAY"� ?c��aS2�e�c���8��BP�MOM�B��@�C�H��Cj��c��3gBT�DUX �2S�_BCKLSH_CS2Fu:��V���C-��esRoz�A�CLA�LMJT@��`� �uC�HKe ����GLRTYpн�8T��5���9_�ùT_UM3��v�C3��1Z���LMT��_LG��%���0�E*�K�=�)�@5F��@8 9�Nb��)hPC��Q)hHТ��5�uC�MC���0�7CN_b��N���;SF�!iV�B��.W���S2�/�ĈCAT�~SH �Å��4 V�q/q/V�0T1��0PA�t�B_P�u�c_f Z�f`�Pe�cݔ�uJG����ѓ�OGއ�TORQU~@�S�i� @e��R� @B�_W u�d�!a��#`��#�`�Ih�Iv�I�#F���S�:��I�0VC"00��֢1ܮ�08��JRKܬ!�,�<�DBXMt�<��M�_DL�!_bGRVg�`��#`��#A��H_%�?��0��CO1S��� ��LN#��� ߥŴ� ��=�������꼰�<�Z���VA�M�YǱ:ȧ��᯻[�T�HET0�UNK2a3�#���#ȰCB��kCB�#Cz�AS��������#����SB8�#��GTSkZAC����&���$DU�phg6�j�(�E�%Q%a_��x�+NEhs1K�t�� y�A}Ŧկ׍�����LPH����^U��Sߥ��������Ҡ�!��(Ʀ�V��V��غ ��V��V��V�
�V�V&�V4�VB�H��������d�����H
�H�H&�H�4�HB�O��O��OTs���O��O��O
�UO�O&�O4�O(ƁF�Ҫ�	���S�PBALANCE�_J�6LE��H_}�SP>!۶^�^>��PFULCb��q���K*1�U�TO_�p�uT1T2�	
22N�q2VP �M�a� i�Z23	q�Tu`O�1Q�IN�SEG2�QREV8�PGQDIF�ep)�1�U�1��`O!BK�qj�w2,�VP��qI�LCHWAR�4B�BAB��u$MECH��J��A��vAX�aPo�����"� � 
�?�1n0UROB�PCRS2X#%Ղ�p�C1_ɒ�T � x ?$WEIGH�@�`#$��\#��I�A�PsIFvA�0LAG�B⎂S�B:�BBILƕ%OD�`�Ps"STD0s"P:�pt  � (N�C!L �P 
P2<�Aɑ  2��Tx&/DEBU�#L|0�"=5�MMY9C59qN��$4�`$D|1� a$0ېl�   �DO_:0AK!� <_ �&� H�q�A��B�"� NJS��8_�P�@�#O�p ��� %�T�7P?Q�TL4F0TgICK�#�T1N0%�3=p�0N�P� u3�PR\p�A��5��5�U0PROMP�CE~�� $IR"��A�p8BX`wBMAI�F��A�BQE_� �OCX�a�@RU�CO�D�#FU�@�&ID�_�P�E82B> G_�SUFF�� h�#�AXA�2DO�70/�5� �6GR�#� �DC�D��E��E-���DU4� �_ H_�FI�!9GSOR�D�! R 236�s�HR�AN0$ZD�T�E'�8�!X5��4 *WL_N�A�1�0�R�5DEF_I�X�RF�T�5�"��6�$�6�S�5�UFISm�#�m1|��40c�3�T6�44􁆂�"�D� ?rfd�#D�O|@ l2LOCKE����C�?OG2a�B�@UM�E�R�D�S�D�U�D >b�B�c�E�S�Dd�B �&2v2a�C�ʑ�E�R��E�S�C9wwu�H�0P@} d�0,a��F0W�h��u�c���T�E�qY4� >�!LOMB_�r�w�0s"VIS��IT�Ys"AۑO�#A_�FRI��~SI,a�n�R�07��07�)3�#s"W�W�Q���%�_���AEAS {#�B��|�x`WB8��45�55�6|#OR�MULA_I����G�W� h �
>75COEFF�_O�1&)��1��Gdo�{#S� 52CA� �:?L3�!GRm� ?� � $�`�v2X�0TM�g���e��2�c��3ERIT��d�T� �  �L�L�Dp`S��_SVLkd��$�v� �.����� � ��SE;TU,cMEAG@�@�Πt �!HRL � �3 (�  0��@l��l��aw��R�0$�a�a}d]�d��B��Ay`Gax`��[�:�k@REC[Qq�=R0MSK_A y��� P_!1_USER�����*���VEL�����-�!��IzP� �M�T�1CFG��� � �0]O�NGOREJ �0l���~[�� 4 e�8��"�XYZ<S��� 3����_ERRK!� U ѐ�1�@Ac�Ȱ�!�>�B0BUFINDX���R0� MORy�� H_ CUȱ�1���dAyQ?�I>Q	$ +�a����� �\�G{�� � $SI�h��@2	��VOv�q�- OBJyE| w�ADJUF2�yĈ�AY�����D��OUKP����AMR=�T��-���X2DIR����X8f�1  DYNt�0�-�T� ��R��0� ~���OPWOR��� �,B0SY�SBU����SOP�o���z�Uy�XP�`K���PA�q��Ӭ���OP�@U����}�"1��IMA�G۱_ �п"IM�.���IN������RGOVRD"ё�	���P����  >gplcC��L�`BŰ?l�PMC_E�P�1EN��Mr�1212�R�"�SL| ��� ��R OVSL=S��rDEX\a`��2�:�_"���P#����P������2�C� �P>���#�_Z�ERl���:����� @��:��O�PR	Iy��
[�g@e����s�P�PL���  $FREEY�EEU�=!Z��L����T�� ATU9Sk�,1C_T�����B������p�Vc18��P��� Dc1������LQ����MQ��ۡL�XE��x�5I�P�W�` ��UP��H`&aPX;@���43�� �PG�Y��g�$SUB����q���JMP�WAIT~ ���L�OW���1wē CV!F_A�0��R�Z��CC �R$��28IGNR_PL��/DBTB� P*a�#BW@.t�U�0-�IG��!@I�TNLN,�RBѡb�yN!@��PEED~ >��HADOW� ��t���E������PwSPD��� L_ �A�нP���	#UN�q � �RP (�L�YwPa���qPH�_PK���b�RE�TRIE��x������H�0NFI���� ���V �$ 2}�d�DBGLV<?LOGSIZz�baKKTU���$D�n�_TXV�EM�!Cڡ��� �-R�#�r>��CHECKz��(�L���ϰq)ҹL��NPA�`T0J"������IP����
�AR�"�BC =S�a��O�@����ATTS�u䡳&� w�^a��3-#UX^�4�fP9L�@Z�� $d��q?SWITCH�h��W��AS������4LLB���� $BA�Dvc��BAMi��6I��(@J5��N�UB�6[F
A_KNOWhK3qB"�U��AD+H�c� D��IPAYGLOAq�9p�C_����GrѼGZ�CLqA�j��PLCL_6� !4��BOA?�T*7�VFYCӐ�J(p��D�I�HRՐ�G$�TB��6�J(�zQ�_J�A �B�AND����T�BQ����PL@AL_ ���0 =�TAe��pCꪢD�CE���J3ܭP�V� T�PDcCK^�)b��COM��_ALPH�ScBaE<�߁�_�\�X�|x\� � ����OD_1�J2�DDM�AR<�h�e�f�c^Q�TIA4�i5�i6��MOM(��c�c��c�c�cV�B� AD��cv�cv�cPUB�P�R�d<u�c<u�b%�8�3���� L$PI$��pc���G�y��I�yI�{I�{I�s�`�A���v��v�J�b��a��HIG�3��� 0���5�0�f�?��5N�5�SAMP D Ƣ�0����;@�S ��с6���1� ��� ���`���`1�@K�P��`腽P�H��IN1��P��8�T��/��:�z�Q�z���G�AMM&�S���$GET�����D�^d>�
$�PIBRt��I��$HI��!_���1��E=��1A�9�*�LW�W� N�9�{�*�Zb���QCdCHK0�j�ݠnI_��M�JļR oh�Q ��sJ�-v㩾�S �$�X �1�N�I�RC�H_D$RN���^�LE��i��p�Zh8�ţMSW�FL/M�PSCRF�75�Ҽ ��3�" Ķ�6��`��ع�����0SV��Pp'������GRO�g�S_SA=AH�=��NO^`Ci�_d =��no�O�O�x�ʚ�`�p�B�u�ȐcDO�A��!�ں�*�tҀ:�Z1f�;�7����C ��LO�nt� � �YL�snQ ��� ���"��<s�	�����nQ૰<N3M_Wl�����\p��(�o�MC��P���Q����rhpM.�pr� ��!ȅ�$�WM��ANGL�!�AM�6dK�=d@K�DdK��TT7�Nk@P��3�#�PXC OEc¼QZ��hp	nt� -���OM���� �ϣϵ����`� c�Z0�0hp^a_�2� | a�J��i���c���c J��j�����jA�s�(�{���s��@{��P�1�PMON_�QU�� � 8�60QCOU��Q�THxHO��B H�YS�0ESPBB U�E- 3�f0O�4� � c P�^�RUoN_TO��	o ��� P�@���INDE�#_PG�RA���0��2��N�E_NO��ITxf��o INFO���a"�����H�O�I� (*�SLEQ!�*�*����OS��l4� 4�60ENABy� PTION�3��r���^GCF�!� �@60J�Q���R�d!��u�P�EDIT�� ��� ��KAQ"� �E�(�NU'(AUT<Y�%COPYAQ�(2,�qe�M�N< @+^��PRUTm� C"�N�OU�2$G���$
�RGADJZ��u2X_��IX�P���&���&W�(P�(�~��&9�� 
�N�P_�CYCy�e1RG�NSc�{�s�LG�O£�NYQ_FREQSrW@��X1�4�L�@�2P0�!�c@�"�CRE��Mà�IF�q�NA���%�4_Gf�STA�TU~�f��MAI�L��|CIq�=LA�ST�1a*4ELE�Mg� ��QrFEASIt;�ւΰ ��B"�F�AF����I� ��O2Z�E u�&vBAB��PE� =��VA�FzQ�I��TqU�[��R��S�FRMS_TRpC�Qc���C��Z�
��1�D X� ,2ns؆�	MB? 2� `��� N�3V�R2WR*����p�R^W�wj�DOU�2^�N�,2PR`�h=�1GRID��oBARS!�TYu$Z�Op��j�} E_�4!� �R�TO��>d� � �����POR�c~vbS�RV�0)"dfDI[�T�`;aNd�pXg
��Xg4Vi��Xg6Vi7�Vi8:av�Fʒg�~z $VALU�C�0�3Dr�ad��C !pf���S�1�-ȆAN/��b�1R��]11ATOTALX����=sPWE3I�Q>StREGENQzfr��X�H�]5	v( cTR�CS�Qq_S3��wfp�V�!��r��BE�3�PG0B�( nsV_H�PDA(��p�S_Ya���i6�S��AR(�2� }�"IG_SE�3ȿpb�5_� �tC_��V$CMPl��D�Ep�G���IšZ�~�X�
��Fm�HA{NC.� p Q�r�2���INT�9`cq�F���MAsSK�3�@OVRMP �PD�1-��W�QaХT�l�_RF�{>�V�PSLGP�g�9�j5��,�;p�DpS���4��U���.�}�TE���`�#��`k���J^�Y�y3IL_Mx4�s��p��TQ( ���@ԍ���V.�C<�P_h �R�F�M]�V1\��V1j�2y�2j�3*y�3j�4y�4j����p۲������ܲIN�VIB8�6�#�T�*�2&�22�3&�32�4&�42��6����SJ�  �T ?$MC_FK `� �L>�J�х1p�Mj�Iу��zS ���1���KEEP�_HNADD��!H鴓@�C��0	��Q����
�O!�v ঱�p
�և
�REM!�	�Cq�RF�]�b��U�4e	�HPWD�  �SBM����PCOLLAB�*�p��/q�2I�T/0��Q"NO1�F�CALp⎵��� �, �FLv�A$�SYN���M��C�k��RpUP_DL�Y��zDELAh9�Dq�2Y AD(�}��QSKIPO�� �`� O��N1T����c�P_� � �׾ ��cp���q�ٞ ��o`��|`�ډ`�ږ`��ڣ`�ڰ`��9�!��J2R0  �lX�@TR3H��1AH� ��H���PRDC\q��� � R�R, 5��R�1��E��5TRGE�_C�㎃RFLG"���W��5TSPC�1U�M_H��2TH2�N}Q�;� 1� �;��Q02 � D� ˈ�鞗@2_PC3W�S����1Y0L10_C�w2��,��� �� $\� U@��V 7�����0���  c�\����� rd��CG�+��7���DZ Gs�RUVL1b[�1h���10]�_DS�������PK ;11�� lڰ�0���q��AT?��$ �Q[7�� ��K 5Tx���HOME�S *�c2h�n`����� _3h���!3�E ��c4h��hz���� y�b5h���	/�/-/?/ N`6h�b/t/�/�/�/�/
�7h��/�/??L'?9? ���!8h�\?n?�?�?�?�?W�S����  ��Aa{p�����_�Ed� T=�nD4v&nCIO䑎II@`�O��_OP�E�C.r���WPOWE	��� X@�f�_�$$Cd�S����j@��3�f3� �@�SI���GP0�~QIRTUAL�O�
QAAVM_WR�K 2 7U� 0  G�5Qn_zXk_.�] �\	�P�]�_3�8P��_�_�Ve�\#m/o�Q5ojo|ōdHPBS�� 1�Y� <Xo�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q���@������˯ݯ�bC$ЯAXLM�@खn�c  d�IN��s�	��PRE
��E�J�-�_UP��[�7QHPIOC�NV_����	�P�r�US>��g�cIO�)�V 1U[P $E`��Qս9lҿ8P?�� �����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�m��LARMRECOV a�$�-����LMDG �ɰ�LM_IF ���ை ����zv����%�6�, 
  6�_��r漅�������̍$w���׏��8��J�\�n����NGT�OL  a� 	? A   ��ț��PPINFO ={ <v���8�1�$�  I�3� a�"rP���t���������ί���>�o�� ��j�|�������Ŀֿ������0�B�PzP�PLICATIO�N ?����+�Ha�ndlingTo�ol �� 
V�9.30P/04�ǐM�
8834�0�å�F0����2�02�ťʚϬ�7�DF3��M̎�No�neM�FRA�M� 6��Z�_�ACTIVE�b � sï�  p�U_TOMODz�A����m�CHGAPO�NL�� ��OUPLED 1ey� ������g��CUREQ 1	�e{  T����	p��w���#rw����e�HN���{�H�TTHKY��$r��\[�m����O�	� '�-�?�Q�c�u����� ��������#) ;M_q���� ��%7I [m���/� ��/!/3/E/W/i/ {/�/�/�/?�/�/�/ ??/?A?S?e?w?�? �?�?O�?�?�?OO +O=OOOaOsO�O�O�O _�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_oo#o5oGoYo ko}o�o�o�o�o�o�o 1CUgy �������	���-�?�Q�c���1�T�O��|�p�DO_CLEAN��n���NM  �� �B�T�f�x���%�DSPDRYR��&m�HI���@/��� ��,�>�P�b�t����������ίj�MAX@a�ۄ�������Xۄ�������p�PLUG�G��܇�ӌ�PRC*��B� ��ׯ�F�OK���ȔSEGF��K�������.������,�>�v���LAPӟ澨�Ϥ϶� ���������"�4�F��X�j߯�TOTAL��7���USENU
Ӱ�� ���ߖ�1��RGDISPMM�C����C����@I@Ȓ��Oѐ������_STRING� 1
��
�kM��Sl�
A�_ITEM1K�  nl�g�y���� ��������	��-�?��Q�c�u����������I/O SIG�NALE�Tr�yout Mod�eL�Inp��S�imulated�P�Out�OVERRА =� 100O�In� cyclP��Prog Abo�rP���Sta�tusN�	Hea�rtbeatJ�MH Faul��Aler�	��� ���*<N` ׃G�ׁY� c�����// //A/S/e/w/�/�/�/�/�/�/�/wWOR ��G�-1�?U?g?y? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O�NPOE��@E; �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_�oo&o8oJo�BDEV�Nu`�Obo�o�o�o �o�o�o,>P bt������>�PALT�� E?�A�S�e�w����� ����я�����+��=�O�a�s����GRI�G뽑1������ 	��-�?�Q�c�u��� ������ϯ����)�����R�a�՟;� ��������ѿ���� �+�=�O�a�sυϗ��ϻ���O�PREG ��y���-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�����$ARG_-0D ?	�������  �	$��	[���]��������S�BN_CONFIQG��� ���CII_SAVE  ��)����TCELLSET�UP ��%  OME_IO�����%MOV_H8n�����REPd������UTOBACK�Y���#�FRwA:\�� ��,��)�'`l ��&�� 7"� �24/07/�25 10:26:54�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� ,,		�����O�G�O __#_%_7_q_[_�_ _�_�_�_�_�_�_%o����D�@TSK � �M&,O��UP3DT�@EGd�`�F�XWZD_ENB8ED��fSTADE��ܖe��XIS�UNOT 2��&�(�� 	\o��; &_J�n���\��dMETc�2LfE� P�!��E���ySCRDCFG� 1�� �A�&�:�����@ԏ�����Q=� ��H�Z�l�~�����	� Ɵ-����� �2�D�0��域���GR�`�`X�O���0NA����s	��_EDC@�1n�� 
 ��%-�0EDT-`q����%�p��(��-��������������  ��B��2����*�?"� D���*�q���ϧ���3bϮ�@Ͻϯd?���@��=�O���sϏ�4.� ��{�����W���	����?ߏ�5��j�G�� ��#������}�6��6��Z�����Z� ���I��7��� ��&��λ�&m�������8^ҿ���� �͇�9K�o��!9*�w����S���;��CR ����B/T//�/���w//��РNO_�DEL����GE_�UNUSE���I�GALLOW 1���   (�*SYSTEM�*)�	$SER�V_GR�;B0�@REGK5$m3)�B0�NUMp:�3�=P�MU� )�LA�Y�p)�PM�PALD@�5CYC10�.�>�0�>CULSU�?�=�2�A�M3LOWDBOX�ORIt5CUR_�D@�=PMCNV6�6D@10�>�@T4DLI�`=O_9�	*PROGRA�J4PG_MI�>�OPAL�E_U�PB7_B>$F�LUI_RESU`�7p_z?�_�TMRY>h0�,�/�b�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv����������"LAL_OUT 1;�l���WD_ABO�R�0?d�ITR_�RTN  �����g�NONSTO�Ǡ�� 8CE_�RIA_I0���ۀ��ŀFCFG ��۔��o_LIMY22ګ� �  � 	i�J��<e�g��5�� 9���������
���u��P}AQPGP 1�����Q�c�u�b4�CK0����C1���9��@���PC��CUV��]��d��l��as��P���C[٤Um��v�������_�� C����-�m��?�ÂHE� �ONFI�Pq�G�G�_P�@1� �%�������ǿٿ�����G�KPAU�SaA1�ۃ  �2�W��Eσ�iϓ� �ϟ����������#߀I�/�m��eߣ��M~��NFO 1"�;�� �7��������/�A8�Δ�e���8�Ώ8m��� �DC@8D���DH  �3�G�´-�?�ŀO��c�COL_LECT_�"�[�����EN�@��y�ܮ�k�NDE���"�3�"1234567890� �\1�� ��֕@�(��)M�r�\,L�^��� ]+������������C  2�Vhz� �����
c .@R�v��������� |����IO !����q���u/�/�/�/�C'TR�2"'-(�׀^)
��.R�#�R-�*W� 9_MOR�$� �;�l5�� l9�?r?�?�?�?�;E2T��%S=,W�?@��@��C׀K)Dց
C�R�&u�XOWAWB_C4  A&��׀�x׀A"@Cz + B�@C@�B8��A�C  @&���׀ց:d�43? <#�
�E��P�I�O�C=AI��'GM�?�C�(S=���Qd�=AT_DEFPR/OG �;%�/m_|APINUSE��V�ۅ�TKEY_TOBL  s�ہ����	
�� �!"#$%&'()*+,-./��:;<=>?@A�BCDPGHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������Ga���͓���������������������������������耇���������������������!�PLCK�\���P΋PSTAn��T_A�UTO_DO��NFsIND���n���R_T1wT2�N����5ŀTRL^CPLETE���z�_SCREEN ��kcs�cÂU��MMEN�U 1)O� < �[_#�q��,�a��� >�d���t���ӏ���� 	�����Q�(�:��� ^�p�������̟�ܟ �;��$�q�H�Z��� �������Ưد%��� �4�m�D�V���z��� ٿ��¿�!���
�W� .�@ύ�d�vϜ��Ϭ� �������A��*�P� ��`�r߿ߖߨ����� ���=��&�s�J�\� �����������'��,�p_MANUAL�EqDB
12�v��iDBG_ERR�LIP*�{h! �0�������g�N_UMLIM�s:Q�OE�@DBPXWO_RK 1+�{���>Pbt��-DBwTB_�q ,���kC3!VD!DB__AWAYo�h!oGCP OB=��A�_AL���o�k�Y�p�uO@`�_�� +1-�+@
-k�-6[��_M+pI�S�`�@"@�ON�TIM�w�ODɼ�&
�U;MO�TNEND�_:R�ECORD 13��{ ��[CG�O�f!T/[K��/�/ �/�/_(�/�/f/?�/ ??Q?c?�/?�??�? ,?�?�?OO�?;O�? _O�?�O�O�O�O(O�O LO_pO%_7_I_[_�O _�O�__�_�_�_�_ l_!o�_,o�_io{o�o �oo�o2o�oVo /A�oeP^�
 ���R���=� �a�s��������*� ߏN���'���ԏ]� ̏��������ɟ۟v� ��n�#���G�Y�k�}����TOLERE�NC�B�0� L���g�CSS_C�NSTCY 24J	�t���.�� ����0�>�P�b�x� ��������ο�����(�:�äDEVI�CE 25ӫ ��ϟϱ������π����/�AߟģHNDGD 6ӫ�� CzT�.!ơLS 27t�S����߀������/�U�ŢPARAM 8G�b�A�Ք�RBTw 2:8��<���CkA�� ·�  �� A���.S�B���A�B�  ���������.��  ����A�A�C����c�u�l���C�A�D�(�k�pz�A�A��HA�c��A�	�? (uL^p��|�A�Bt/�D���C��_ 	 �A=��ABffA#33AҊ���A�A�C%f��a��A�J���7B]��B��BffBᴠ�33C$.@R� (����A� ����
/��// )/;/�/_/q/�/�/�/ �/�/�/�/<??%?r? I?[?m??�?�?�?�? �?&O8O�PObOMO�O qO�O�O�O�O�O_� OOL_#_5_�_Y_k_ �_�_�_�_ o�_�_6o ooloCoUogo�o�o �o�o�o�o �o	 h�O�w���� �
��.�	__I'� 1_�q��������ˏ ݏ���%�r�I�[� ���������ǟٟ&� ���\�3�E�W���� ȯ���ׯ�"��F� 1�j�E�s�����m��� ����ѿ�0���f� =�O�a�sυϗ��ϻ� �������'�9�K� ��o߁�����[���� (��L�7�p��m�� ������������$��� ��l�C�U���y��� �������� ��	V -?�cu��� �
��@+dO �s������� �*///`/7/I/[/ m//�/�/�/�/?�/ �/?!?3?E?�?i?{? �?�?�?�?�?�?�?FO �jOUOgO�O�O�O�O �O�O__�'O9OO =_O_�_s_�_�_�_�_ �_�_�_oPo'o9o�o ]ooo�o�o�o�o�o �o:#5��O� ���� ��$���H�Fz�$DCSS�_SLAVE �;���w���`�_4D � w���AR_M�ENU <w�  >�؏���� �2�^r�Ǐ\�n�\���SH�OW 2=w� � fr[q����Ə �����,�>�D�b�t��� ����ҟϯ� ���)�P�M�_�q� ��������˿ݿ�� �:�7�I�[ς�|Ϧ� �ϵ���������$�!� 3�E�l�fߐύߟ߱� ���������/�V� P�z�w������� ������@�:�d�a� s�����������\��� *�H�N�K]o� �������2 8�GYk}�� ����"�1/ C/U/g/y/�/��/�/ �/��//?-???Q? c?u?�/�?�?�?�/�? ?OO)O;OMO_O�? �O�O�O�?�O�?�O_ _%_7_I_pOm__�_ �O�_�O�_�_�_o!o 3oZ_Woio{o�_�o�_ �o�o�o�oDo- Se�o��o��� ���.�=�O����CFG >������q��dM�C:\��L%04�d.CSV\��pc��������A ՃCH݀z�v�w�#�_  ����:�J�8�S���JP�j�)���p7�-��n�RC_OUT [?z������a�_C_FSI �?�� |�����@�;� M�_���������Я˯ ݯ���%�7�`�[� m��������ǿ�� ���8�3�E�Wπ�{� �ϟ����������� �/�X�S�e�wߠߛ� �߿��������0�+� =�O�x�s������ �������'�P�K� ]�o������������� ����(#5Gpk }����� � HCUg�� ������ // -/?/h/c/u/�/�/�/ �/�/�/�/??@?;? M?_?�?�?�?�?�?�? �?�?OO%O7O`O[O mOO�O�O�O�O�O�O �O_8_3_E_W_�_{_ �_�_�_�_�_�_oo o/oXoSoeowo�o�o �o�o�o�o�o0+ =Oxs���� �����'�P�K� ]�o�����������ۏ ���(�#�5�G�p�k� }�������şן ��� ��H�C�U�g����� ����دӯ��� �� -�?�h�c�u������� ��Ͽ�����@�;� M�_ψσϕϧ����� ������%�7�`�[� m�ߨߣߵ������� ���8�3�E�W��{� ������������� �/�X�S�e�w����� ����������0+ =Oxs���� ��'PK ]o������ ��(/#/5/G/p/k/ }/�/�/�/�/�/ ?�/�??H?C?U3�$D�CS_C_FSO ?����1� P [?U?�?�?�?�?�? O
OO.OWOROdOvO �O�O�O�O�O�O�O_ /_*_<_N_w_r_�_�_ �_�_�_�_ooo&o OoJo\ono�o�o�o�o �o�o�o�o'"4F oj|����� ����G�B�T�f� ��������׏ҏ��� ��,�>�g�b�t��� ������Ο����� ?�:�L�^����������ϯʯܯg?C_RPI~>�?�;�d�_� 
�}?.�p����ݿj>SL�@���9�b� ]�oρϪϥϷ����� �����:�5�G�Y߂� }ߏߡ���������� ��1�Z�U�g�y�� �����������	�2� -�?�Q�z�u������� ������
)R M_q����� ��*%7Ir m�����/ �ϛ�,�/W/�/{/ �/�/�/�/�/�/?? ?/?X?S?e?w?�?�? �?�?�?�?�?O0O+O =OOOxOsO�O�O�O�O �O�O___'_P_K_ ]_o_�_�_�_�_�_�_ �_�_(o#o5oGopoko }o�o�o�o�o�o �o HCUg�� ������ �����NOCODE �@������PRE_CHKg B��3�A 3���< ��7��������� 	 <�����?#ۏ%�7� �[�m�G�Y������� ٟ�ş�!����W� i�C�����y�ïկˏ ������A�S�-�_� ��c�u���ѿ����� ��=��)�sυ�_� �ϻϕ��������'� 9���E�o�I�[ߥ߷� ����������#���� Y�k�E���{���� ��������C�U�� =�����w��������� 	����?Q+u� a������ );_qg�Y� �S����%/� /[/m/G/�/�/}/�/ �/�/�/?!?�/E?W? 1?c?�?���?�?o? �?O�?�?AOSO-OwO �OcO�O�O�O�O�O_ �O+_=__I_s_M___ �_�_�_�_�_�?�_'o 9oo]oooIo�o�oo �o�o�o�o#�oG Y3E��{�� ���o�C�U�� y���e����������� 	��-�?��K�u�O� a���������͟�� )��1�_�q��}��� ����ݯ�ɯ�%��� 1�[�5�G�����}�ǿ ٿ�������E�W� 1�{ύ�G�u����ϯ� �����/�A��-�w� ��c߭߿ߙ������� ��+�=��a�s�M�� ��ϑ�������'� �3�]�7�I������ ������������G Y3}�i���� ����C/ y�e����� ��-/?//c/u/O/ �/�/�/�/�/�/�/? )?�?_?q?K?�?�? �?�?�?�?�?O%O�? IO[O5OO�OkO}O�O �O�O�O_�O3_E_;? -_{_�_'_�_�_�_�_ �_�_�_/oAooeowo Qo�o�o�o�o�o�o�o +7aW_i_� �C�����'� �K�]�7�i���m�� ɏۏ�������G� !�3�}���i���ş ������1�C��g� y�S�e���������� ѯ�-���c�u�O� ������Ͽ�ןɿ� )�ÿM�_�9�kϕ�o� �����Ϸ������ I�#�5�ߑ�kߵ��� ��������3�E��� Q�{�U�g������� �����/�	��e�w� Q��������������� +Oa�I� ������ K]7��m� ����/�5/G/ !/k/}/se/�/�/_/ �/�/�/?1???g? y?S?�?�?�?�?�?�? �?O-OOQOcO=OoO �O�/�/�O�O{O�O_ �O_M___9_�_�_o_ �_�_�_�_oo�_7o Io#oUooYoko�o�o �o�o�o�O�o3E i{U����� ���/�	�S�e�?� Q�������я㏽�� ��O�a������� q���͟������� 9�K�%�W���[�m��� ɯ�����ٯ�5�+� =�k�}���������� ���տ�1��=�g� A�Sϝϯω����Ͽ��������Q�c�����$DCS_SG�N CS������g�29�-JUL-24 ?09:35 EӘ�}5��10:30������� X�S��������������Д���ÿ������ � {�VERSIO�N ��V�4.2.10�E�FLOGIC 1�DS��  	D���X�k��X�z�M�PROG_�ENB  ���b��Л�ULSE � ���M�_A�CCLIM��������WRS�TJNT����w�EMO���ѷ�L���INIT E�Z�O��OPT_�SL ?	S�1�
� 	R575��Ӆ�74��6��7R��5A��1��2���l���G�h�TO  �t���.H�V?�DKEX��d����FPATH A�ڇA\4���H�CP_CLNTI�D ?+�b� �l�����IAG_GRP 2JS�� ����[�D� � D�� D  B�  B�@gff��/B�@�[��W�@�q���B�N�C��-Bz��Bp�@e`��m�p3m7 7890123456��*�[��  A�o�mAj1A�dA]�
A�W|�AP�A�J-AC/A;�A4H���_@�  A��A�YA3!_A�@@v��B4�� ���t���
�uƨA�pffAj�yA�eK�A_�A�Y��AS� MC��AF��A@ �O�+/=/O$O�c K��w(@�X?8�?�@��y�/�/p�/�/�/8�;d�2��5?@~ff@�x1'@q��@�kC�@d�D@]��@Vv�6?�H?Z?l?~?8s�0l���@e@^���@W\)@O���@H�0?<@7?K�@.V�?�?��?�?
O8S@�M00G<@A��@�<1@5��@�/l�@(Ĝ@!�0�\NO`OrO �O�Ox'g�L_K�;_�_ �__g_�_�_�_�_o �_�_�_YokoIo�o�o+o�oX�"� 2�1x7A�@J>��R
q�?�33?Y���r��J7'���2q63p4�F�>r��LJ@�p��Zr�
=@��@�Q�jq��@VG Ah�@��@�T�= c<��]�>*�H>V�>�3�>���~J<���<�p�q�x��� �?�� �C�  <(��U�� 4Vr��33��@
���A@��?R�oD��mR�x� ��Q��t����Z�Џ���؏�,��i?�7>N�>�(�>�@Z��=���J��G�v�G�J�B�E������a��@ǐ@����@��@Q�?�L ���ŲI@�P���&���'��@�K����Ag�q��PC�  C�̇�Cuy�
���ʯ  ?����	��Գ�4���X��v���+�� A�¿�������π@�+�F��Iϗ�C�T_CONFIG� K3����eg��ST�BF_TTS��
@����"�������{��MAU���MS�W_CF��L � �OCVIE�W	�MI�U�� 㯛߭߿��������� ���0�B�T�f�x�� ������������� ,�>�P�b�t������ ����������(: L^p���� �� �6HZ l~�����X�/��RCB�N��!��F/{/j/�/��/�/�/�/��SBL�_FAULT �O9*^�1GPMS�K��7��TDIAOG P��U�����qUD1�: 6789012345q2�q���%P�ϭ?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O �a6�I'��
�?_��TREC	PJ?\:
j4\_�7_[ �?�_�_�_�_�_�_o o(o:oLo^opo�o�o��o�o�O�O_ _�U�MP_OPTIO1N��>qTRB���:9;uPME��.�Y_TEMP  È�3B����p�A�pytUNI�'��ŏq6�YN_B�RK Qt�_�EDITOR q&qh��r_2PENT 1�R9)  ,& �/0��d�[�`�J��� n��������ȏ�� )�;�"�_�F�����|� ����ݟğ֟���7� �F�m�T���x���ǯ ���ү�!��E�,��i�P��pMGDI_STA�u~��q���p�NC_INFO �1SI��b��������Կⷮ���1TI� ��o#��0�
0�d�o}Ϗϡϳ� ����������1�C� U�g�yߋߝ߯����� ����Hu� �2�D�R� j�R�x�������� ������,�>�P�b� t�������������Z� �#5Ga�k} ������� 1CUgy�� ������	//-/ ?/Yc/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? ��?O%O7OQ/GOmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�?Ooo /o�_[Oeowo�o�o�o �o�o�o�o+= Oas����� �_�_��'�9�So]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�K�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�C�5� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ�������� �!�;�M�W�i�{�� ������������� /�A�S�e�w������� ��������+E� Oas����� ��'9K] o����1��� �/#/=G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?��?�?	OO5/ ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�?�_ �_oo-O#oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���_�_���� 7oA�S�e�w������� ��я�����+�=� O�a�s��������� ߟ���/�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������͟׿���� '�1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߫�ſ ���������;�M� _�q��������� ����%�7�I�[�m� ������߯������� �)�3EWi{� ������ /ASew���� �����/!+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?/��?�?�? �?/#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �?�_�_�_�_Oo-o ?oQocouo�o�o�o�o �o�o�o);M _q���_��� �	o�%�7�I�[�m� �������Ǐُ��� �!�3�E�W�i�{��� ��ß՟矝��� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}� �ߩ����������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u����߫��� ��������);M _q������ �%7I[m �������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?���? �?�?�?�OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�?�?�_�_�_�_�? �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�_� ����_�	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q��y�����˟� ۟��%�7�I�[�m� �������ǯٯ�����!�3�E�W�i��� ��$ENETMO�DE 1U��  ���������»��R�ROR_PROG %��%������TABLE  ���Q�c�uσ���SEV_NUM� ��  �������_AUT�O_ENB  �̵��ݴ_NO�� �V������ W *���������	�����+���(�:ߞ��FLTR����H�IS�Ð�����_A�LM 1W�� e����̍�+;߀��������0�?�_\����  �����²u꒰TCP_V_ER !��!���@�$EXTLOGo_REQv�������SIZ����ST�K�������T�OL  ��Dz�~��A ��_BWDU�*�Z�V�ǲ?�DID� X��Z�����[�ST�EPl�~�����OP�_DO���FAC�TORY_TUN�v�d��DR_GR�P 1Y��`�d �	p�.° �*�u���RH�B ��2 ���� �e9 ���bt�o�� �����J�5nY@��oA�@��@D�v@��`�u
 E�����uȸo���_/�(/(B� � F!A���33�R"�33-@UU�Tn*@� /ȷ>�u.�>*��<���ǆ-�F@� �"�5W�%�-J���NJk�I�'PKHu��IP�sF!���-�?�?�/9�<�9�89�6C'6<,�5���/  �������D��� f������FEATUROE Z�V�Ʊ�Handl�ingTool ��5��Engl�ish Dict�ionary�74�D St�0ard��6�5Analog� I/O�7�7gle Shift O�uto Soft�ware Upd�ate%Imati�c Backup��9SAground� Edit�0�7C_amera�0F�?�CnrRndIm�XC�Lommon �calib UI�C�FnqA�@Monoitor�Ktr�0?Reliab@�8�DHCP�IZat�a Acquis��CYiagnos�OA�1[ocume�nt Viewe��BWual Ch�eck Safe�ty�A�6hanc�ed�F�:�UsnPF�r�@�7xt. D7IO �@fiRT�Wwend�PErr�@QLQR�]�Ws�Yr�0��P E�:FCTN_ Menu�Pv S�8gTP In'`f�acNe�5GigE�`nrej@p Mas_k Exc�Pg�W�HT^`Proxy� SvoT�figh�-Spe�PSki�D�eJP�Pmmun�icN@ons�hu�rE`'`_�1abconnect 2x�ncr``struH�2z>peeQPJQU��4KAREL C�md. L�`ua��husRun-Ti��PEnvkx(`el� +R@sP@S/W��7License��Sn\�PBook(System)�:MACROs,�b?/Offse@�uaH�P8@_�pMR�@��BP^MechSt�op�at.p6R�ui�RKj�x�P�0P@)��od@witchȘ�>�EQ.���Op�tmЏ>��`fil�n\=�gw�uult�i-T�`tC�9PC�M funHwF�o�3T�R?�f�Regi��pr�`I�rigPF�V����0Num S�elb����P Ad�ju�`���J�t�atu��
�iZ�5R�DM Robot>�0scove�1F��ea7��PFreq� Anly�gRe�m`��Qn�7F�R�S�ervo�P���8S�NPX b�rNSN^`ClifQɮB�Libr�3鯢0 �q�����o�ptE`sGsag?��4�� -C���;��/I_mB�M�ILIBk�E�P OFirm6BU�PEc�Acck@sKTPT9X_C�eln����F��1�V�orqu>@imula�A�A�u��Pa�qU�j@t�Ã&�`ev.B��.@riP޿USB port �@�iP�PagP��R �EVNT�ϗ�nexcept�P��t�X�ſX�]VC�Ar�b�bf�V2PҦ�$�����SܠSCصV�S�GEk�a�UI�;Web Pl!��ާ���Խ`�TeQfZD?T Appl�d�:x�ƺ� �GridV�play�R�WD4�R
�.�:n�EQ+��r�-10iA/7L�*��1Graphi�c���5dv�SDC�SJ�ck�q�5la�rm Cause�/��ed�8Asc�ii�a��Load�nP�Upl,�Ol�0�AGu�6N�`���yFyc@�r�����P�V��Jo��m� c��R���c���m�./������Q�2*u:eRA`J��P�ٶ4eqinL�����8NRT��9O}n�0e Hel�H�J�`oI�allet�iz?�H�����_�t�r�[ROS Eth�q��T@e�ׅ�!��n�%�2D�tPkgp&Upg~��(2DV-�3D� Tri-jQEA�ưDef.qEBa)pdei��� �b�ImπF�f��n�sp.q=�464M?B DRAMZ,#�FRO5/@ell��<�Mshf!r/�'c�%3@pLƖ,ty�@s˒xG��m��. [�� ��BU���Q�B�=mai�P߫�]hQ����@q6wlu��H��^`�xR�?eL� Sup������0�P�`cr��@�R���b�x���pr1uest�Crt~QQ��ߋL!��4O��q$�K��l� Bui7�n��A'PLCOO�EVl%��sCGU�OCRG�Ob��DR��O
TLS_&��BU/_��K�qN_&d�TA�OxVB�_�Wp�ܑZ���_TCB�_ �V�_�W���WF+o�V��O�W._�W�ņoTE�H�o�f�O�gt�oT	Ej�xVF�_w�_xV�GoTwBTw~oxVH�xVIA��v�xVLN�yUMz�boH�f_xVN�xVP�H��^xVR&xVS��܇ʏ��W��v���gVGF:�L�P2_�h��h�V�h��_g�D���h�FFoh��g�R�D�� TUT��0�1:�L�2V�L�TB�GG��v�rain�UI��
%HMI���pon��m��f�"�F�&K�AREL9� �TPj��<5�
"E�<�N� {�r���������̿޿ ���A�8�J�w�n� �ϭϤ϶�������� �=�4�F�s�j�|ߩ� �߲���������9� 0�B�o�f�x���� ���������5�,�>� k�b�t����������� ����1(:g^ p�������  -$6cZl� �������)/  /2/_/V/h/�/�/�/ �/�/�/�/�/%??.? [?R?d?�?�?�?�?�? �?�?�?!OO*OWONO `O�O�O�O�O�O�O�O �O__&_S_J_\_�_ �_�_�_�_�_�_�_o o"oOoFoXo�o|o�o �o�o�o�o�o KBT�x��� ������G�>� P�}�t�������׏Ώ �����C�:�L�y� p�������ӟʟܟ	�  ��?�6�H�u�l�~� ����ϯƯد���� ;�2�D�q�h�z����� ˿¿Կ���
�7�.� @�m�d�vψϚ��Ͼ� �������3�*�<�i� `�r߄ߖ��ߺ����� ���/�&�8�e�\�n� ������������� +�"�4�a�X�j�|��� ������������' 0]Tfx��� ����#,Y Pbt����� ��//(/U/L/^/ p/�/�/�/�/�/�/�/ ??$?Q?H?Z?l?~? �?�?�?�?�?�?OO  OMODOVOhOzO�O�O �O�O�O�O_
__I_ @_R_d_v_�_�_�_�_ �_�_oooEo<oNo `oro�o�o�o�o�o�o A8J\n �������� �=�4�F�X�j����� ��͏ď֏����9� 0�B�T�f�������ɟ ��ҟ�����5�,�>� P�b�������ů��ί ����1�(�:�L�^����   �H552}���21n��R78��50���J614��ATU]PͶ545͸6���VCAM��CRIn�UIFͷ28	ƷNRE��52��R�63��SCH��DwOCV]�CSU���869ͷ0ضEI�OC9�4��R69���ESET���J�7��R68��MA{SK��PRXY!�]7��OCO��3�h����̸3�J6˸�53��H2�LCH^��OPLG�0֯MHCR��S{�MkCS�0��55ض�MDSW���OP��MPR�M�@�0n̶PCM �R0���ض��@�51�5u1<�0�PRS�ǻ69�FRD�FwREQ��MCN��{93̶SNBAE�^3�SHLB��M��tM���2̶HTC��TMIL����TP�A��TPTX��EL��Ѐ�8������wJ95,�TUT׻95�UEV��U�EC��UFR�V�CC��O��VIP��CSC,�CSGt8�r�I��WEB�7HTT�R6C�N��CGIG��IP�GS)RC�DG��H77��6ضR�85��R66�Ru7��R:�R530�K680�2�q�J��*H�6<�6,�RJح�j0�4�6o64\��5�NVD��R6��R84Tg�����8�90\���J9&3�91� 7+����,�D0oF�CL9I���CMS�� n�STY��TO䶴q���7�NN�O�RS��J% ��j�O]L(END��L���Sf(FVR��V3�D���PBV,�A�PL��APV�C�CG�CCR|�C�D��CDL@CS�Bt�CSK��CT�CTBL9��U0,(�C��y0L8C��TC� �y0�'TC(7TC���CTE\��07T�Eh��0��TFd8FJ,(GL8GI�8H�8�I��E@�87�CTM�,(M�8M@8N�8P�HHPL8Rd8(TSrd8W�I@VGF�GP2��P2���@�H�{7VPD�HF �V�PSGVPR�&VT���YP��VTB7Vs�IH��VI aH'VK��V���_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U?�g?y?�9  H55hT�1�1[Un�3R78�<50�9�J614�9ATU\�T�4545�<6�9�VCA�D�3CRIf,KUI8T�528-J�NRE�:52JR�63�;SCH�9D�OCV�JCU�48�69�;0�:EIOt�TsE4�:R69J�ESET�;KJ7�KR68�JMAS�K�9PRXYML7.�:OCO\3�<�J�)P�<3|ZJ6�<5u3�JH�\LCH\Z�OPLG�;0�ZM�HCR]ZSkMC�S�<0,[55�:MgDSW}k�[OP�[GMPR�Z�@�\0�:7PCMLJR0�k)P��:)`�[51K51�|0JPRS[6�9|ZFRD<JFR�EQ�:MCN�:9=3�:SNBA}K�[/SHLB�zM�{�@�ll2�:HTC�:T�MIL�<�JTPA��JTPTX�EL��z)`�K8�;�0�JJ�95\JTUT�[9�5|ZUEVZUE�C\ZUFR<JVCuC��O<jVIP,�wCSC\�CSGlJ��@I�9WEB�:H�TT�:R6{L��C�G{�IG[�IPGmS��RC,�DG�[�H77�<6�:R8�5�JR66JR7�[R|R53{6%8|2�Z�@Jml,|6|6\JR�\	P|�4L�6�64��5n�kNVDZR6+k�R84<���IP,�8f��90���KJ9�\91��̫7[KIP\J�D0�F��CLI�lKCMS�J9��:7STY,�TO�:�@��K7�LNN|ZOR�S<jJ��MZZ|OL�K�END�:L�S��FVR�JV3D�,�KKPBV\�AP�L�JAPV�ZCC�G�:CCRjCD��CDL̚CSBn�JCSK�jCTK��CTB��\���\�Ch�z���CL�TCLJl�l�TC��TCZ�CTE�J��|�TEX�J��<�TF��F\̥G��G��l�Hl�Ip�z)�l�k�CTM\�UM\�M��Nl�P,�eP��R��;�TS�ܹW��̚VGF��P2��P2�z ��VPDFLJVPn;�VPR��VT�;\� �JVTB��V�K�IH�VِM�<�VK,�V{��8#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew ������� +=Oas�� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G?�Y?k?}?�5�0�STD�4LANG�4�9�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~��������� �2�D�V�RB=T�6OPTNm�� ������Ǐُ���� !�3�E�W�i�{�����8��ß�5DPN�4� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳ڈ8�� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s���������pͯ߯��  ���*�<�N�`�r���9�9���$FEAT�_ADD ?	��������  	��ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu�����DEMO Z��?   ���} ��'��0�]�T�f� �������������� #��,�Y�P�b����� ������������ (�U�L�^��������� ���ܯ���$�Q� H�Z���~�������� ؿ��� �M�D�V� ��zόϦϰ������� �
��I�@�R��v� �ߢ߬��������� �E�<�N�{�r��� �����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo~o �o�o�o�o�o�o�o! *WN`z�� �������&� S�J�\�v��������� �ڏ���"�O�F� X�r�|�������ߟ֟ ����K�B�T�n� x�������ۯү�� ��G�>�P�j�t��� ����׿ο���� C�:�L�f�pϝϔϦ� ������	� ��?�6� H�b�lߙߐߢ����� ������;�2�D�^� h����������� ��
�7�.�@�Z�d��� �������������� 3*<V`��� �����/& 8R\����� ����+/"/4/N/ X/�/|/�/�/�/�/�/ �/�/'??0?J?T?�? x?�?�?�?�?�?�?�? #OO,OFOPO}OtO�O �O�O�O�O�O�O__ (_B_L_y_p_�_�_�_ �_�_�_�_oo$o>o Houolo~o�o�o�o�o �o�o :Dq hz������ �
��6�@�m�d�v� ������ُЏ��� �2�<�i�`�r����� ��՟̟ޟ���.� 8�e�\�n�������ѯ ȯگ����*�4�a� X�j�������ͿĿֿ ����&�0�]�T�f� �ϊϜ����������� �"�,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/
??A? 8?J?w?n?�?�?�?�? �?�?�?OO=O4OFO sOjO|O�O�O�O�O�O �O__9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿����&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t����������   ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�����y  �x�q��� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p��P����q�p�x ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p���������������$F�EAT_DEMO�IN  ��� �����IND�EX���I�LECOMP �[���B���8 SETU�P2 \B~L�  N w�5_AP2BCK� 1]B	  #�)����%����E �	���5 �Y�f��B ��x/�1/C/� g/��/�/,/�/P/�/ t/�/?�/??�/c?u? ?�?(?�?�?^?�?�? O)O�?MO�?qO O~O �O6O�OZO�O_�O%_ �OI_[_�O__�_�_ D_�_h_�_�_
o3o�_ Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0����ׯQ	� P� 2>� *.VRޯ(���*+�Q���W�{��e��PC������OFR6:��ؾg�����T   �2�����\� ��d�*.F��ϕ�	ó����qo�ߓ�STM� 9���ư%�d��ψ���HU߻�Jש�f�x���GIF�A�L��-����ߑ��JPG ����Lձ�n�����#JS�H�����6����%
JavaS�criptt���C�Se���Kֹ�v� %�Cascadi�ng Style Sheets���j�
ARGNAMOE.DT'��OЁ\;��[�k|(>k DISP*rU�Oп��� �
�TPEINS.X3ML/�:\C�cCustom Toolbar���	PASSWOR�D���FRS:�\�� %Pa�ssword Config/c�Q/ �J/�/���/:/�/�/ p/?�/)?;?�/_?�/ �??$?�?H?�?l?�? O�?7O�?[OmO�?�O  O�O�OVO�OzO_�O �OE_�Oi_�Ob_�_._ �_R_�_�_�_o�_Ao So�_woo�o*o<o�o `o�o�o�o+�oO�o s��8��n ��'���]���� �z���F�ۏj���� ��5�ďY�k������ ��B�T��x����� C�ҟg�������,��� P���������?�ί �u����(���Ͽ^� 󿂿�)ϸ�M�ܿq� ��ϧ�6���Z�l�� ��%ߴ��[����� �ߵ�D���h����� 3���W����ߍ��� @����v����/�A� ��e������*���N� ��r�����=��6 s�&��\� �'�K�o� �4�X��� #/�G/Y/�}//�/ �/B/�/f/�/�/�/1? �/U?�/N?�??�?>? �?�?t?	O�?-O?O�?�cO�?�OO(O�O�F��$FILE_DG�BCK 1]����@��� < �)
S�UMMARY.DyG�OsLMD:�O�;_@Diag� Summary�<_IJ
CONSLOG1__&Q_�_NQ�Console� log�_HK	T�PACCN�_o%�o?oJUTP A�ccountin��_IJFR6:I�PKDMP.ZI	PsowH
�o�oKU[`�Exceptio�n�oyk'PMEMCHECK5o�_*_K��QMemory� DataL�F�/l�)6qRIP�E�_$6�Zs%��q Packe�t L�_�DL�$y�	r�qSTAT����S� %~�rStatusT��	FTP���:����Vw�Qmmen�t TBD؏� �>I)ETHERNE���
q�[��NQEthern��p�Pfigura��oODDCSVRAF̏��ďݟd���� verify �all��{D�.���DIFF՟��͟xb��s��diffd���
q��CHG01 Y�@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ��VTRNDIAG.LS�̿޿s�^q=3� Ope���q� SQnostic�EWY�)VD;EV7�DATt�Q�xc�u�g�Vis��?Device�Ϫ�IMG7ºo����y�z�s�Imag�n��UP��ES��~T�FRS:\��� �OQUpdates List ��IJg�FLEXEVENQ�X�j߃�f��F� UIF E�v���B,�s��)
PSRBWLOD.CM��sL�������PPS_RO�BOWEL��GL�o�GRAPHIC�S4Dy�b�t���%4D Gra�phics Fi�leu��AOɿ��rGIG���u�
>YvGigE�ة�~�BN�? )��HADOW������\sShadow Chang���vbQRCMERR�n�\s�� CFG Er�ror�tail�� MA��C?MSGLIB� �"^o� ���T�)�ZD�����/XwZD�6 ad�HPNOTI���
/�/Zu�Notific8��H/��AGUO�/ yO?�O'?P?OOt?? �?�?9?�?]?�?O�? (O�?LO^O�?�OO�O 5O�O�OkO _�O$_6_ �OZ_�O~_�__�_C_ �_�_y_o�_2o�_?o ho�_�oo�o�oQo�o uo
�o@�odv �)�M��� ��<�N��r���� ��7�̏[������&� ��J�ُW������3� ȟڟi�����"�4�ß X��|������A�֯ e�����0���T�f� ���������O��s� �ϩ�>�Ϳb��o� ��'ϼ�K����ρ�� ��:�L���p��ϔߦ� 5���Y���}���$�� H���l�~���1��� ��g���� �2���V� ��z�	�����?���c� ��
��.��Rd�� ���M�q �<�`��� %�I��/� 8/J/�n/��/!/�/ �/W/�/{/?"?�/F? �/j?|??�?/?�?�?��$FILE_F�RSPRT  ����0�����8MDON�LY 1]�5�0� 
 �)M�D:_VDAEX?TP.ZZZ�?�?�_OnK6%N�O Back f�ile 9O�4S�6Pe?�OOO�O�?�O __?>_�Ob_t__�_ '_�_�_]_�_�_o(o �_Lo�_po�_}o�o5o �oYo�o �o$�oH Z�o~��C� g��	�2��V�� z������?�ԏ�u��
���.�@��4VIS�BCKHA&C*�.VDA�����F�R:\Z�ION\�DATA\v�����Vision VD�B��ŏ��� '�5��Y��j���� ��B�ׯ�x����1� ��үg�������X��� P��t���Ϫ�?�ο c�u�ϙ�(Ͻ�L�^� �ς��)���M���q�  ߂ߧ�6���Z���� ��%��I�������:�LUI_CONF�IG ^�5|m��� $ h� �3��������/�A�D$ |xq�s��� ��������a���  $6��Gl~�� �K��� 2 �Vhz���G ���
//./�R/ d/v/�/�/�/C/�/�/ �/??*?�/N?`?r? �?�?�???�?�?�?O O&O�?JO\OnO�O�O )O�O�O�O�O�O_�O 4_F_X_j_|_�_%_�_ �_�_�_�_o�_0oBo Tofoxo�o!o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� �����ʏ܏��� $�6�H�Z�l������ ��Ɵ؟ꟁ�� �2� D�V�h���������¯ ԯ�}�
��.�@�R� d�����������п� y���*�<�N�`��� �ϖϨϺ�����u�� �&�8�J���[߀ߒ� �߶���_������"� 4�F���j�|���� ��[�������0�B� ��f�x���������W� ����,>��b t����O���(:�  �xFS�$FL�UI_DATA �_������uRESULT 2`��� �T��b����/"/ 4/F/X/j/|/�/�/� ��/�/�/�/?"?4? F?X?j?|?�?�?�?�=}?� 0�� ��?�;��O-O?O QOcOuO�O�O�O�O�O �O�O�#
O_/_A_S_ e_w_�_�_�_�_�_�_�_���?g�?;o �?boto�o�o�o�o�o �o�o(:L]o p�������  ��$�6�H�oi�+o ��Oo��Ə؏����  �2�D�V�h�z����� ]ԟ���
��.� @�R�d�v�����Y��� }�߯�����*�<�N� `�r���������̿޿ 𿯟�&�8�J�\�n� �ϒϤ϶������ϫ� �ϯ1�C��j�|ߎ� �߲����������� 0�B��f�x���� ����������,�>� ��G�!�k���W߼��� ����(:L^ p��S����  $6HZl~ �O���s�����/  /2/D/V/h/z/�/�/ �/�/�/�/�
??.? @?R?d?v?�?�?�?�? �?�?����9O� `OrO�O�O�O�O�O�O �O__&_8_�/\_n_ �_�_�_�_�_�_�_�_ o"o4oFoOO)O�o MO�o�o�o�o�o 0BTfx�I_� ������,�>� P�b�t�����Woio{o ݏ�o��(�:�L�^� p���������ʟܟ� ��$�6�H�Z�l�~� ������Ưدꯩ�� ͏/��V�h�z����� ��¿Կ���
��.� @�Q�d�vψϚϬϾ� ��������*�<��� ]����C��ߺ����� ����&�8�J�\�n� ���Q϶��������� �"�4�F�X�j�|��� M߯�q����ߗ� 0BTfx��� �����,> Pbt����� ���/��%/7/�^/ p/�/�/�/�/�/�/�/  ??$?6?�Z?l?~? �?�?�?�?�?�?�?O  O2O�;//_O�OK/ �O�O�O�O�O
__._ @_R_d_v_�_G?�_�_ �_�_�_oo*o<oNo `oro�oCO�OgO�o�o �O&8J\n �������_� �"�4�F�X�j�|��� ����ď֏�o�o�o�o -��oT�f�x������� ��ҟ�����,�� P�b�t���������ί ����(�:���� ��A�����ʿܿ�  ��$�6�H�Z�l�~� =��ϴ����������  �2�D�V�h�zߌ�K� ]�o��ߓ���
��.� @�R�d�v����� �������*�<�N� `�r������������� ������#��J\n �������� "4EXj|� ������// 0/��Q/u/7�/�/ �/�/�/�/??,?>? P?b?t?�?E�?�?�? �?�?OO(O:OLO^O pO�OA/�Oe/�O�/�O  __$_6_H_Z_l_~_ �_�_�_�_�_�?�_o  o2oDoVohozo�o�o �o�o�o�O�o�O+ �_Rdv���� �����*��_N� `�r���������̏ޏ ����&��o/	S� }�?����ȟڟ��� �"�4�F�X�j�|�;� ����į֯����� 0�B�T�f�x�7���[� ��Ͽ������,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸��߉��� ����!��H�Z�l�~� �������������  ���D�V�h�z����� ����������
. �����s5��� ���*<N `r1������ �//&/8/J/\/n/ �/?Qc�/��/�/ ?"?4?F?X?j?|?�? �?�?�?��?�?OO 0OBOTOfOxO�O�O�O �O�O�/�O�/_�/>_ P_b_t_�_�_�_�_�_ �_�_oo(o9_Lo^o po�o�o�o�o�o�o�o  $�OE_i+_ ��������  �2�D�V�h�z�9o�� ��ԏ���
��.� @�R�d�v�5��Y�� }�����*�<�N� `�r���������̯�� ���&�8�J�\�n� ��������ȿ��鿫� ���F�X�j�|ώ� �ϲ����������� ݯB�T�f�xߊߜ߮� ����������ٿ#� ��G�q�3Ϙ����� ������(�:�L�^� p�/ߔ�����������  $6HZl+� u�O������  2DVhz�� ������
//./ @/R/d/v/�/�/�/�/ }���?�<?N? `?r?�?�?�?�?�?�? �?OO�8OJO\OnO �O�O�O�O�O�O�O�O _"_�/�/?g_)?�_ �_�_�_�_�_�_oo 0oBoTofo%O�o�o�o �o�o�o�o,> Pbt3_E_W_�{_ ����(�:�L�^� p���������woɏ�  ��$�6�H�Z�l�~� ������Ɵ�矩� �2�D�V�h�z����� ��¯ԯ���
��-� @�R�d�v��������� п�����ן9��� ]���ϖϨϺ����� ����&�8�J�\�n� -��ߤ߶��������� �"�4�F�X�j�)ϋ� Mϯ�q�s������� 0�B�T�f�x������� �������,> Pbt����{� �����:L^ p�������  //��6/H/Z/l/~/ �/�/�/�/�/�/�/? ��;?e?'�?�? �?�?�?�?�?
OO.O @OROdO#/�O�O�O�O �O�O�O__*_<_N_ `_?i?C?�_�_y?�_ �_oo&o8oJo\ono �o�o�o�ouO�o�o�o "4FXj|� ��q_�_�_�_	��_ 0�B�T�f�x������� ��ҏ�����o,�>� P�b�t���������Ο ��������[� ���������ʯܯ�  ��$�6�H�Z��~� ������ƿؿ����  �2�D�V�h�'�9�K� ��o�������
��.� @�R�d�v߈ߚ߬�k� ��������*�<�N� `�r�����y��� ������&�8�J�\�n� ���������������� !�4FXj|� �������� -��Q�x��� ����//,/>/ P/b/!�/�/�/�/�/ �/�/??(?:?L?^? ?A�?eg?�?�?  OO$O6OHOZOlO~O �O�O�Os/�O�O�O_  _2_D_V_h_z_�_�_ �_o?�_�?�_o�O.o @oRodovo�o�o�o�o �o�o�o�O*<N `r������ ���_o�_/�Y�o ��������ȏڏ��� �"�4�F�X�|��� ����ğ֟����� 0�B�T��]�7����� m�ү�����,�>� P�b�t�������i�ο ����(�:�L�^� pςϔϦ�e�w����� �Ͽ�$�6�H�Z�l�~� �ߢߴ��������߻�  �2�D�V�h�z��� ����������
����� ��O��v��������� ������*<N �r������ �&8J\� -�?��c����� /"/4/F/X/j/|/�/ �/_�/�/�/�/?? 0?B?T?f?x?�?�?�? m�?��?�O,O>O PObOtO�O�O�O�O�O �O�O_O(_:_L_^_ p_�_�_�_�_�_�_�_  o�?!o�?EoOlo~o �o�o�o�o�o�o�o  2DV_z�� �����
��.� @�R�os�5o��Yo[� Џ����*�<�N� `�r�������g̟ޟ ���&�8�J�\�n� ������c�ů����� ��"�4�F�X�j�|��� ����Ŀֿ������ 0�B�T�f�xϊϜϮ� �������ϵ���ٯ#� M��t߆ߘߪ߼��� ������(�:�L�� p�����������  ��$�6�H��Q�+� u���a���������  2DVhz�� ]�����
. @Rdv��Y�k� }������/*/</N/ `/r/�/�/�/�/�/�/ �/�?&?8?J?\?n? �?�?�?�?�?�?�?�? ���CO/jO|O�O �O�O�O�O�O�O__ 0_B_?f_x_�_�_�_ �_�_�_�_oo,o>o PoO!O3O�oWO�o�o �o�o(:L^ p��S_����  ��$�6�H�Z�l�~� ����aoÏ�o珩o�  �2�D�V�h�z����� ��ԟ���	��.� @�R�d�v��������� Я������׏9��� `�r���������̿޿ ���&�8�J�	�n� �ϒϤ϶��������� �"�4�F��g�)��� M�O����������� 0�B�T�f�x���[� ����������,�>� P�b�t�����W߹�{� ������(:L^ p������� ��$6HZl~ ���������� ��/A/h/z/�/�/ �/�/�/�/�/
??.? @?�d?v?�?�?�?�? �?�?�?OO*O<O� E//iO�OU/�O�O�O �O__&_8_J_\_n_ �_�_Q?�_�_�_�_�_ o"o4oFoXojo|o�o MO_OqO�O�o�O 0BTfx��� ����_��,�>� P�b�t���������Ώ ���o�o�o7��o^� p���������ʟܟ�  ��$�6��Z�l�~� ������Ưد����  �2�D���'���K� ��¿Կ���
��.� @�R�d�vψ�G��Ͼ� ��������*�<�N� `�r߄ߖ�U���y��� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������	�� -��Tfx��� ����,> ��bt����� ��//(/:/��[/ /AC/�/�/�/�/  ??$?6?H?Z?l?~? �?O�?�?�?�?�?O  O2ODOVOhOzO�OK/ �Oo/�O�O�?
__._ @_R_d_v_�_�_�_�_ �_�_�?oo*o<oNo `oro�o�o�o�o�o�o �O�O�O5�O\n �������� �"�4��_X�j�|��� ����ď֏����� 0��o9]���I�� ��ҟ�����,�>� P�b�t���E�����ί ����(�:�L�^� p���A�S�e�w�ٿ��  ��$�6�H�Z�l�~� �Ϣϴ����ϗ����  �2�D�V�h�zߌߞ� �������ߥ���ɿ+� �R�d�v����� ��������*���N� `�r������������� ��&8��	�� }?������ "4FXj|;� ������// 0/B/T/f/x/�/I�/ m�/��/??,?>? P?b?t?�?�?�?�?�? �?�/OO(O:OLO^O pO�O�O�O�O�O�O�/ �O�/!_�/H_Z_l_~_ �_�_�_�_�_�_�_o  o2o�?Vohozo�o�o �o�o�o�o�o
. �OO_s5_7�� �����*�<�N� `�r���Co����̏ޏ ����&�8�J�\�n� ��?��cşן���� �"�4�F�X�j�|��� ����į֯������ 0�B�T�f�x������� ��ҿ��۟����)�� P�b�tφϘϪϼ��� ������(��L�^� p߂ߔߦ߸�������  ��$��-��Q�{� =Ϣ�����������  �2�D�V�h�z�9ߞ� ����������
. @Rdv5�G�Y�k� ����*<N `r������� �//&/8/J/\/n/ �/�/�/�/�/�/�� �?�F?X?j?|?�? �?�?�?�?�?�?OO �BOTOfOxO�O�O�O �O�O�O�O__,_�/ �/?q_3?�_�_�_�_ �_�_oo(o:oLo^o po/O�o�o�o�o�o�o  $6HZl~ =_�a_��_���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П����<�N� `�r���������̯ޯ ���&��J�\�n� ��������ȿڿ��� �"��C��g�)�+� �ϲ����������� 0�B�T�f�x�7��߮� ����������,�>� P�b�t�3ϕ�WϹ��� ������(�:�L�^� p���������������  $6HZl~ ���������� ��DVhz�� �����
//�� @/R/d/v/�/�/�/�/ �/�/�/??�!� E?o?1�?�?�?�?�? �?OO&O8OJO\OnO -/�O�O�O�O�O�O�O _"_4_F_X_j_)?;? M?_?�_�?�_�_oo 0oBoTofoxo�o�o�o �oO�o�o,> Pbt����� �_�_�_��_:�L�^� p���������ʏ܏�  ���o6�H�Z�l�~� ������Ɵ؟����  ����e�'����� ��¯ԯ���
��.� @�R�d�#�u������� п�����*�<�N� `�r�1���U���y��� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ���������	��� 0�B�T�f�x������� ����������> Pbt����� ����7��[ �������  //$/6/H/Z/l/+ �/�/�/�/�/�/�/?  ?2?D?V?h?'�?K �?�?�/�?�?
OO.O @OROdOvO�O�O�O�O }/�O�O__*_<_N_ `_r_�_�_�_�_y?�? �?�_o�?8oJo\ono �o�o�o�o�o�o�o�o �O4FXj|� ��������_ o�_9�c�%o������ ��ҏ�����,�>� P�b�!��������Ο �����(�:�L�^� �/�A�S���w�ܯ�  ��$�6�H�Z�l�~� ������s�ؿ����  �2�D�V�h�zόϞ� ���ρ������ɯ.� @�R�d�v߈ߚ߬߾� �������ſ*�<�N� `�r��������� ����������Y�� ���������������� "4FX�i� ������ 0BTf%��I�� m����//,/>/ P/b/t/�/�/�/�/� �/�/??(?:?L?^? p?�?�?�?�?w�?� �?�$O6OHOZOlO~O �O�O�O�O�O�O�O_ �/2_D_V_h_z_�_�_ �_�_�_�_�_
o�?+o �?OoOo�o�o�o�o �o�o�o*<N `_������ ���&�8�J�\�o }�?o����wڏ��� �"�4�F�X�j�|��� ����q֟����� 0�B�T�f�x������� m�����ۯ�Ǐ,�>� P�b�t���������ο ���ß(�:�L�^� pςϔϦϸ�������  ߿�	��-�W��~� �ߢߴ����������  �2�D�V��z��� ����������
��.� @�R��#�5�Gߩ�k� ������*<N `r���g��� �&8J\n ����u������ ��"/4/F/X/j/|/�/ �/�/�/�/�/�/�? 0?B?T?f?x?�?�?�? �?�?�?�?O��� MO/tO�O�O�O�O�O �O�O__(_:_L_? ]_�_�_�_�_�_�_�_  oo$o6oHoZoO{o =O�oaO�o�o�o�o  2DVhz�� ��o���
��.� @�R�d�v�������ko ͏�o�o�*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� ����C���|��� ����Ŀֿ����� 0�B�T��xϊϜϮ� ����������,�>� P��q�3��ߧ�k��� ������(�:�L�^� p����e�������  ��$�6�H�Z�l�~� ����a߫߅�������  2DVhz�� �������. @Rdv���� ���������!/K/ r/�/�/�/�/�/�/ �/??&?8?J?	n? �?�?�?�?�?�?�?�? O"O4OFO//)/;/ �O_/�O�O�O�O__ 0_B_T_f_x_�_�_[? �_�_�_�_oo,o>o Poboto�o�o�oiO{O �O�o�O(:L^ p������� �_�$�6�H�Z�l�~� ������Ə؏����o �o�oA�h�z����� ��ԟ���
��.� @��Q�v��������� Я�����*�<�N���o�1������$F�MR2_GRP �1a���� �C4  �B�[�	 [��߿�ܰE�� Fw@ 5W��S�ܰJ��NJk��I'PKHu���IP�sF!{���?�  W��S�ܰ9�<9��896C�'6<,5�{��A�  ��6��BHٳB�հ��޷�@�33�3�3S�۴��ܰ@UUT'�@��8���W�>u.�>*�߭<����=[��B=���=�|	<�K�<��q�=�mo����8�x	7H�<8�^6�?Hc7��x?��� �������"��F�X����_CFG b»T Q���|��X�NO º/
F0�� ��W��RM_CHKTYP  ��[�ʰ̰܂���ROM�_MsIN�[���9�u���X��SSBh��c�� ݶf�[�]����^��TP_DEF_O��[�ʳ��IR�COM���$G�ENOVRD_D�O.�d���THR�.� dd��_E�NB�� ��RA�VC��dO�Z�� ���Fs  G�!� GɃ�I��C�I(i J����+���%������ �QOUU��j¼������<6�i�C`�;]�[�C�հ��հȡ`��[�@ر����.��.R SMT��k_	ΰ�\��$HOST�Ch�1l¹[�̭d� 	�(�+��/Z��/W�e �/??'?9?G:�/j?�|?�?�?�/�?W0	anonymouy  �?�?	OO-O?N�/�/ �/�O�?�/Y?�O�O�O _K?(_:_L_^_p_�O �?�?�_�_�_�_ oGO YOkO}O_lo�O�o�o �o�o�o_�o 2 Dgo�_�_���� �o-o?o�S@��o d�v������o��Џ� ��)�*�qN�`�r� ���������� I�&�8�J�\�n����� ����ȯگ��3�E�"� 4�F�X�j���ß՟�� �ֿ�����0�B� �f�xϊϜϿ���� ������,�s����� ���߽�߿�������� �K�(�:�L�^�p�� ���ϸ������� �G� Y�k�}��l��ߐ��� ��������� 2 U�C��z�����//h!ENT 1m� P!V  7 ?.c &�J�n��� /�)/�M//q/4/ �/X/j/�/�/�/�/? �/7?�/?m?0?�?T? �?x?�?�?�?O�?3O �?WOO{O>O�ObO�O �O�O�O�O_�OA__ e_(_:_�_^_�_�_�_��ZQUICC0 �_�_�_?od1@oo.o�od2�olo~o�o�!ROUTER��o�o�o/!PC�JOG0!�192.168.�0.10	o�SCA�MPRT�\!bpu1yp��vRT�o���� !So�ftware O�perator Panel�mn���NAME !~�
!ROBO��v�S_CFG 1�l�	 ��Auto-st�arted'�FTP2��I�K2� �V�h�z������� ԟ����	���@�R� d�v���	������ �:���)�;�M�_�&� ��������˿�p�� �%�7�I�[��"�4� F�ڿ��������!� 3���W�i�{ߍߟ��� D���������/�v� �Ϛ�w�ߛ��Ͽ��� ������+�=�O�a� ��������������� 8�J�\�n�p�]�� �������� #5X�k}�� ��0/D1/ xU/g/y/�/RH/�/ �/�/�//?�/??Q? c?u?�?���/? �?:/O)O;OMO_O&? �O�O�O�O�O�?pO_ _%_7_I_[_�?�?�? t_�O�_O�_�_o!o 3o�OWoio{o�o�_�o Do�o�o�o����_ERR n���-=vPDUSIZW  �`^�P�Tt�>muWRD ?�΅�Q�  guest�f�������~�S�CDMNGRP �2o΅WpC��Q�`���fKL�� 	P01.0�5 8�Q   ��|��  };|��  z[� ���w����*���Ť�x����[ݏȏ�V�בPԠ���~���)����D�Yr���؊p"�P�l�P���Dx��d�x�*�����%�_GR�OU7�pLyN���	/�o���QUP���UTu� �T�YàL}?pTT�P_AUTH 1�qL{ <!i?Pendan�����o֢!KAR�EL:*�������KC��ɯۯ��V�ISION SET�9����P�>�h� �f����������ҿ�����X�CTRL rL}O�uſa�
�aFFF9�E3-ϝTFRS�:DEFAULT���FANUC� Web Server�ʅ�u�X�� �t@���1�C�U�g��;tWR_CONF�IG s;� ���=qIDL_C_PU_PC���asBȠP�� BH���MIN�܅q��GNR_IOFq{r�`Rx���NPT_SIM�_DO��STAL_SCRN�� �.�INTPM?ODNTOLQ����RTY0����-�N\�ENBQ�-���OLNK 1tL{�p������)�;�|M���MASTE��%���SLAVE �uL|�RAMCOACHEk�c�O^�O_CFG�������UOC�����CMT�_OP���PzY�CL������_AS�G 1v;��q
 O�r����� ��&8J\\W�ENUMzsPy�
��IP����RTRY_CN��M�(=�zs���Tu ������w���p/�p���P_MEMBER�S 2x;�l� $��X"��?�Q'W/�i)��RCA_AC�C 2y�  X�\} j���� 6��"  '
�`�`�&�#�#�/��#�/�$BUF0�01 2z�= �Zu0  uW0Z$:44:4E:4UT:4e:4u:4�:4U�:4�:4�:4�:4��:4�:4�:3[	��4�4)�48�4K��4Z�4k�4{�4���4��4��4��4Ҫ�4�4�4�:3\U*D*D.*D=*DUN*D]*Dn*D}*D��h  hX��:3X�zD�zD�V:3Y�D�D!�DU0�DA�DP�Da�DUq�D��D��D��De��DÒDDY�D%�:4:392$?63 :1@1ERI0ERQ0ERY0 ERa0ERi0ERq0ERy0 ER�0ER�0ER�0ER�0 ER�0ER�0:1�1�R�0 �R�0�R�0�R�0�R�0 �R�0�R�0�R�0�R�0 �R@�R	@�R@�R@ �R!@�R)@:10A5b9@ 5bA@5bI@5bQ@5bY@ 5ba@5bi@5bq@rAxA :1�A�b�@�b�@:1�A �b�@�b�@�b�@�b�@ �b�@�b�@�b�@�b�@ �b�@�b�@�b�@�b�@ �bdQ�bPERP:193-_65GSNrI2WS NrY2gSNri2wSNry2 �SNr�2�SNr�2�SNr �2�S�r�2�S�r�2�S �r�2�S�r�2�S�r�2 c�r	Bc�rB'c�r )B7c>�9BGc>�IBWc >�YBgc>�iBwc��xC �c���B�c���C�c�� �B�c���B�c���B�c ���B�c���B�c���B s��	RsNrR'v��2{�4r�}ŋ���<����o�o��2��HIS!2}� �ܷ! 2024�-07-29�&���П���  8�:` 1;oal�!�3�E�xW�i� 2X�_K��5������Ưد�o�_K���,�>�/� O�!����������ο ����(�_�q�^� pςϔϦϸ�������  �7�I�6�H�Z�l�~� �ߢߴ������!��  �2�D�V�h�z��� ���������
��.� @�R�d�v���k��,P�������������:2L�c�� d� o�dWi{�{���@�����9c�� A.@Rd���� �����//*/ </N/���/�/�/�/ �/�/�/??&?]/o/ \?n?�?�?�?�?�?�? �?�?5?G?4OFOXOjO |O�O�O�O�O�OOO 1O_0_B_T_f_x_�_ �_�_����5p����� o$o6o���w�Aovo �o�o�o��o�o ��`��CUgy ��O�O�o���	� �-�?�Q�c���� ����Ϗ����)� ;�M������������� ˟ݟ���%�\�n� [�m��������ǯٯ ���4�F�3�E�W�i��{�������ÿտ�_I_CFG 2~�[� H
Cycle Time��Busy�I�dl��minz�S�Upƾ�Read(��DowG�C� �W��Count>�	Num ��������`����P�ROG���U��P�)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,1�C�U��g�y�Tä�SDT_�ISOLC  ��Y� ���J2�3_DSP_EN�B  ��T���INC ����c���A   ?�  �=���<#�
|���:�o ��2�D��a/�l���OB���C��O��ֆ�G�_GROUP 1큦�<�*�����t�?�����`Q'�L�^�p�@/����������\��~�G_IN_AU�TO����POSR�E���KANJI_MAS@p2��D�RELMON ��[���by����@����f�Ã�ǉ���d-��K�CL_L NUM���G$KEYLO�GGINGD�P��������LANGU�AGE �U���DEFA�ULT ��QLGf�����S���a}x�  8T�oH  ��`'0����`;�`ߍ�;���
*!(UTg1:\ J/ L/ Y/k/}/�/�/�/�/�/��/�/$>(�H?�VL�N_DISP ����P�&�$�^4OCgTOL�0�aDz�����
�1GBOOK ��d4V�11�07u%O!O3O EOWOiKyM�TËIgF	�5)����O}����2_BUFF ;2��� ��`2O�_�2��6_M�R_ d_�_�_�_�_�_�_�_ �_o3o*o<oNo`o�o��o�o�o���ADCS ������L�O���+=Oa�dI�O 2��k +������� �����*�:�L� ^�r���������ʏ܏����$�6�J�uuE_R_ITM��d�� ����ǟٟ����!� 3�E�W�i�{��������ïկ�����7x�S�EVD��t�TYP����s�������)RSTe�eSC�RN_FL 2�
�}�����/�`A�S�e�wϨ�TP{���b��=NGNA�M��E��dUPS�f0GI��2�����_LOAD��G� %��%RE�QMENU�Ϧ<MAXUALRMb,2�@���
K���'_PR��2  �3�AK�Ci0��qO=_x'X�Ӭ�P 2��;W �*V	����
*����4��*� �'�`�	xN��z�� ����������1�C� &�g�R���n������� ����	��?*c FX������ �;0q\ �������/ �/I/4/m/X/�/�/ �/�/�/�/�/�/!?? E?0?i?{?^?�?�?�? �?�?�?�?OOAOSO�6OwObO�OD�DBG?DEF ��գ���ѤO�@_LDXD�ISA����ssME�MO_AP��E {?��
 �A �H$_6_H_Z_l_~_�_��_K�FRQ_CF�G ����CAM �G@��S�@<�ԃd%�\o�_�P�Ґ�����*Z`/\b **: eb�DXojho�F�o�o �o�o�o�o;�O ��dZ�U�y|��z,(9�Mt��� 1��B�g�N���r��� �����̏	���?�~A�ISC 1���K` ��O�����O����O֟����K�]�_M?STR �3���SCD 1�]� �l��{�����د ïկ���2��V�A� z�e�������Կ���� ���@�+�=�v�a� �υϾϩ�������� �<�'�`�K߄�oߨ� �ߥ��������&�� J�5�Z��k����� ����������F�1� j�U���y��������� ����0T?x6�MK�Q�,��Q��$MLTARM��R�?g� �~s�@���@ME�TPU�@l���4�NDSP_AD�COL�@!CM�NT7 *FN�SW(FSTLI8xi%� �,�����Q��*POS�CF�bPRP�MV�ST51��,� 4�R#�
 g!|qg%w/�'c/�/�/ �/�/�/�/?�/?G? )?;?}?_?q?�?�?�?��?�1*SING_�CHK  {$oMODA�S�e����#EDEV }	�J	MC:WL�HSIZE�Ml ��#ETASK %��J%$123456789 �O�E!GTRIG 1�,� l�Eo#_�y_S_�}�FYP�A�u9D�"CEM_INF� 1�?k`)�AT&FV0E�0X_�])�QE0�V1&A3&B1�&D2&S0&C�1S0=�])A#TZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_ �_�_o�3o��o� ��o��"�4��X� ��ASe֏� ��C�0���f�!� ��q�����s�䟗��� ��͏>��b���s��� K���w���ٯ�ɟ ۟L����#�����Y� ʿ����$�߿H� /�l�~�1���U�g�y� ���ϯ� �2�i�V�	πz�5ߋ߰ߗ���PON�ITOR�G ?�kK   	EOXEC1o�2�3�4�5��@�U7�8�9o� ����(��4�� @��L��X��d��Pp��|��2��2��U2��2��2��2��U2��2��2��2��3��3��3(�#AR�_GRP_SV �1��[ (s��Dq >Nnl���`��Nng5c��v
#A�A_Ds���N��ION_DB�-@�1Ml  ��l QFH" -	e�l 
FH��N BL�"FI-ud1�}E���)PL_NAME !�E�� �!Def�ault Per�sonality� (from FsD)b*RR2��� 1�L�XL��p�X  d��.@Rdv� ������// */</N/`/r/�/�/�/f2)�/�/�/??@,?>?P?b?t?f<�/ �?�?�?�?�?�?
OO@.O@OROdOc	���?"�N
�O�OfP�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_�O �O2oDoVohozo�o�o �o�o�o�o�o
. @o!ov���� �����*�<�N��`�r����� F�s  GT�Gg�Me���ÏՍfd����� (�6������
��n�~�8h����� ���� ��ğ֟�����:����
�]�m�f��	`ট����į��:��oAb	����c? A�  /��� P����r�������^��˿ݿȿ��%��RN�� 1��	X ��, � ���� a� @D�  &t�?�z�`�?f |�fA/��t�{	���;�	l��	 ��xJ������� �� ��<�@���� ���·�K�K ���K=*�J����J���J9��
�ԏC߷��@�t�@{S�\��(Ehє��.���I����>����T;f�ґ��$��3��´  �@��>�Թ�$��  >�����;�U��x`���� �
���Ǌ���� �  {�  @T�����/  �H �l�����-�	'� �� ��I� ��  �<�+�:��È��È=��Q������N �[�?�n @���f����f�k���,�<av�  '��Y����@2��@�0c@�Ш���C��}Cb C��\C�������G�@�~� (lݿ@X*�B�b $/�!��L��Dz�o�ߓ~������( �� -��������!���/��|��恀?�ffG�*<� }�q�"��8����>��bp$��(�(���P��	�������>�?����x�����<
6�b<߈;܍��<�ê<���<�^��I/��A�{��fÌ�,��?fff?_�?&�� T�@�.�"��J<?�\��"N\�3���!��(�|� �/z��/j'��[0?? T???x?c?�?�?�?�?0�?�?3��%F��? 2O�?VO�/wO�)IO�O�EHG@ G@0~��G�� G}� �O�O�O_	_B_-_f_�Q_BL��B[�A w_[_�_b��_�[�_�� mO3o�OZo�_~o�o�o<�o���b��PV( @|po	lo-*cU�ߡA���r5�eCP�Lo�}?����#��3���W�s��6�Cv�q�CH3� j�t�����q�����|^(�hA� �ALf�fA]��?�$��?��;�°�u�æ�)�	�ff��C�#s�
���g\)�"��33C�
�����<�؎�G�B������L�B�s�����	";�H��ۚG��!G���WIYE���C�+�8��I۪I�5��HgMG�3�E��RC�j=�x�
�pI����G��fIV=�?E<YD�C<� ݟȟ����7�"�[� F��j�������ٯį ���!��E�0�i�T� f�����ÿ���ҿ� ���A�,�e�Pω�t� �Ϙ��ϼ������+� �O�:�s�^߃ߩߔ� �߸������ �9�$� 6�o�Z��~����� �������5� �Y�D� }�h����������������
C.(䁳3��/"����u���t��q3ǭ8����q4M�gu���q�Vw�Q�
4p�+4�]$$dR�Pv���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/�/X�/�/�/  %��/ �/+??O?:?s?/�_0�?�?�?�;�?�?@O�? OFO4O�rLO�^O�O�O�O�O�O�J � 2 FsH�GwT�V�M�uaBO�|r�pp�C��S@�R_�poy_�_^_l�_o \!�W�Ƀ�_oo(o�z?_���@@�z�t��p�p�q�p�~
 6o�o�o�o �o�o�o);M�_q�ڊsa �����D��$M�R_CABLE �2�� �]��T�LaMa?��PMaLb�p�Z���&P�C�p�!O4>ÔB]�%���v�l/  ��&P�v�wdN�{0���6��H�XT��6P� C$�Čj�|����t% ��&P��C���=�о�Џ��s9� �T�,�>���b����� ��Ɵ��Ο3�.��P��(�:���^����� �������H�Z��l�*��**} �sOM ��y�����Bj���%% 2345?678901ɿ۵! ƿ���� �� AQ5� �!
�z��not sen�t ���W��TESTFECoSALG� eg;j"AQd��ga%�
���@���$�r�̹�������� 9UD�1:\maint�enances.�xmS�.�@�vj��DEFAUL�T�\�rGRP 2=���  p�Xwk�  �%1st� mechani�cal chec�k��!���������E��Z�(��:�L�^��"��controller�����߰��D�����0 ��$�s�M��L��""8b���v��B�����������/�AC}�a�6����@dv���s�C���ge��. battery�&��E	S(:L^p�	�|�duiz�abl�et  D�а�R���/�"/4/s��gre�as��'f�r#-� |!�/�E��/�/��/�/�/s�
�oi0,�g/y/�/�/t? �?�?�?�?s��
�XֈW��1<X�AO�E
c?8OJO\OnO�OB�t��?O��'O��O_ _2_D_s�O?verhauE��L��R xXЌQ�_���O�_�_�_�_o�X�$�_0o����_o  �_�o�o�o�o�oo�o ?oQocoJ\n� ��o�)�� "�4�F���|��k� �ď֏����[�0� B���f����������� ҟ!���E�W�,�{�P� b�t�����矼��� �A��(�:�L�^��� ��ѯ㯸��ܿ� � �$�s�Hϗ���~�Ϳ �ϴ�������9��]� o�Dߓ�h�zߌߞ߰� ����#�5�G���.�@� R�d�v��ߚ������ ������*�y���`� ��O������������ ?�&u�J��n� ����); _4FXj|�� ��%�//0/ B/�f/���/��/ �/�/�/?W/,?{/�/ b?�/�?�?�?�?�?? �?A?S?(Ow?LO^OpO �O�O�?�OOO+O�O _$_6_H_Z_�O~_�O �O�O�_�_�_�_o o�P�R	 T"oOoao so�_�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z��������ԏ���
�� � ��Q?�  @�a �oW�i��{��fC�����̟�h;*�** �Q�V ��� �2�D��h�z��������_�S� �����կ7�I�[� ����ɯ/���ǿٿ#� ��!�3�}�����{� �ϟ��s�������C� U�g��S�e�w�9ߛߠ�߿�	�߉e�a��$MR_HIST� 2��U�� �
 \jR$ 23�45678901P*�2����)�9c_ ���R��a_����� ����=�O�a��*�x� ����r������� 9��]o&�J� ����#�G��k}4��d�S�KCFMAP  ]�U������`��ON�REL  �����лEXCFENB'
��!�FNC$/$JOG_OVLIM'd�\m �KEY'p%=y%_PAN(�"\�"�RUN`,�+�SFSPDTYPxD(%�SIGN/>$T1MOTb/!��_CE_GRoP 1��U� "�:`��n?�c[?�?�� �?�?~?�?�?�?!O�? EO�?:O{O2O�O�OhO �O�O�O_�O/_�O(_ e__�_�_�_�_v_�_��_�_o�׻QZ_�EDIT4��#T�COM_CFG 1��'%to�o�o� 
Ua_ARC_�!"��O)T_MN�_MODE6�Lj_SPL�o2&U?AP_CPL�o3$�NOCHECK {?� � Rdv���� �����*�<�N��`��NO_WAI�T_L 7Jg50NTF]a���UZ��o_ERR?12���ф��	��-����PR�d����`O����| j�
o��Z9<� �� ?���ϟ����قPARAuMႳ��N����R�=��o��� = e������گ� ȯ��"�4��X�j�F�<�蜿��A�ҿ�"?ODRDSP�c6�/(OFFSET_�CAR@`�o�DI�S��S_A�`A�RK7KiOPEN_FILE4�1�a�Kf�`OPTION�_IO�/�!��M_�PRG %�%c$*����h�WOT�[�E7O��и�Z��  ��� �Z"�÷"�	� �W"�Z����RG_DSBOL  ��ˊ����RIENTT5O ZC����A �U�`IM_ED���O��V�?LCT ���Gb�ԛa�Zd��_P�EX�`7�*�RAT��g d/%*��UOP ���{��������������$�PAL�������_?POS_CHU�7�����2>3�L��XL�p��$�ÿU�g�y����� ����������	- ?Qcu����Y2C���"4 FXj|��� ��� //$/6/H/ Z/l/~/�Y���.��/�/ςP�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO�/�/ LO^OpO�O�O�O�O�O �O�O __$_6_H_Z_ )O;O�_�_�_�_�_�_ �_o o2oDoVohozo`�o�o�_<���o�m ���~B Pw�m�m���~�jw8��w����� �2�T��p��w���H��t	`���̏ޏ��:�o����� �|2���A�  I� �j�`�������� �џ���@��#��)�Or�1��_�� 8���, �\Ԡ��� @D�  ��?����~�?� ���!D�������G�  �;�	l��	 ��xJ�젌����� �+<� ���%�	��2�H(��H3k�7HSM5G�2�2G���GNɁ3%�R��oR�d�2�C%f��a��{�ׄ���|��/��3��¸��4��>���К������3�A�q½{{q�!ª��ֱ� "�(«�=�2�ܤ��� ��{ � @�Њ���  ��Њ�2����.�	'� � ���I� � � �V�,�=�������˖ß��� � �y��n �@"��]�<߭˄�ȅ���-�N�Д�  �'�Ь�w�ӰC��C��\C߰��Ϲ�x�ߤ!���@�4�� (l0�_@X+�B��@B�I�;�)�j客z+����쿱����������( �� -��#������&�!�]�9��  q�?�ffaH�Z���� ��������8� ����>�|P��}�	(� ��P�������\�?��� x�� ���<
6b<�߈;܍�<��ê<���<G�^�*�gv�A)�ƙ�脣��F�?f7ff?}�?&� ���@�.��J<�?�\��N\� �)���������� �ޤy�N9r] �������/ &/�J/5/n/�	�g/�/c(G@ G�@0i�G�� G}���/??<?'?`?�K?�?o?BLi�B��A�?y?�?|��?K �?ů�/QO�/xO�?�O�O�O�Om��b��n�t @|�O'_�O@K_6_H_�_lS��A��RS�i�Cn_�_j_0O�]?��ooAol,où�Wi���To3C���`CHQo>J�d�`a�a@I�ܚ>(hA� ��ALffA]���?�$�?����ź°u�æ��)�	ff��?C�#�
�op�g\)��33C��
�����<���nG�B����L�B��s�����	0źH�ۚG���!G��WI�YE���C��+�½I۪�I�5�HgM�G�3E��R�C�j=�~
�p�I���G��f�IV=�E<YD�#Zo���
� �U�@�y�d������� ��я�����?�*� c�N���r�������� ̟��)��9�_�J� ��n�����˯���گ �%��I�4�m�X��� |���ǿ���ֿ��� 3��W�B�Tύ�xϱ� ����������	�/�� S�>�w�bߛ߆߿ߪ� ��������=�(�a�:L�(q��)�����Z��x����a3�8���<���a4Mgu�����a�VwQ�(�4p�+4�]B� B���p����������U%PbP���QO%�x�1[FjR��������  C���I4m X�8
O������.//>/d/R/�Rj/|/�/�/�/��/�/:  2 {Fs�gGT�&6�M�eBmp�R�P�aC��3@�_p?�?@�?�?�?�?�=�S��OO)O;OMO�c?̯��@@�j�R�`�`�1�`�^
 TO�O�O�O�O �O_#_5_G_Y_k_}_p�_�_�j�A ������D��$PA�RAM_MENU� ?B���  DEFPULSE�[�	WAITTM�OUTkRCV�o SHEL�L_WRK.$CUR_STYL`;DlOPTZ1Zo�PTBooibC?oR?_DECSN`�� �l�o�o�o& OJ\n�������QSSREL_�ID  >�
1���uUSE_PRO/G %�Z%�@��sCCR` �
1�S�S�_HOST �!�Z!X���M�T  _���x������>L�_TIMEb ��h��PGDEBU�G�p�[�sGINP?_FLMSK�E�qT� V�G�PGAr�e 5��?��CHS�^D�TYPE�\�0��
�3�.�@�R� {�v�����ï��Я� ���*�S�N�`�r� ���������޿�� +�&�8�J�s�nπϒ����G�WORD ?�	�[
 	PyR2��MAI�`ΓSU�a��TE�Ԁ���	Sd�CCOL��C߸�L�� C�~�h�d�*�TRACECToL 1�B��QW ��0'��|�Ӂ�DT Q�B���М�D � �������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OE��.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�"Op� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r����������� ��&�8�J�\�n��� �������������� "4FXj|�d� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o��c�$PGTRA�CELEN  ��a  ����`��f_UP ����q�'pq   p�a_�CFG �u�	s�a p�Lt��ceqxc}  ��qu4rDEFSP/D �?|�ap���`H_CON?FIG �usW �`�`d�tM��b �a�qP�t�cq��`��`IN~7pTRL �?}�_q8�u�PE�u��w�qLt�q\qv�`LID8s�?}�	v�LLB 1¾�y ��B��pB4Ńqv ��އ؏	�s <�<0p  ?� �'���A�o�U�w� ������۟��ӟ��#�	�+�Y�v�񂍯�� ��ï
��������/�~u�GRP 1ƪ���a@�j���hs�aA�
�D�� D@� �Cŀ @�٭�^�t������q�p����.� ���Ⱦ´���ʻB�)�	����?�)�c��a>��>�,��Ϻ������ =49X=H�9��
����@�+� d�O���s߬�o߼�����  Dz���`
��8���H�n�Y�� }�������������@4��X�C�|���)���
V7.10b�eta1Xv �A������!������?!G�>¿�\=y�#��{�33A!��@���͵��8wA���@� A�"s�@Ls���� ��"�4FXLsAp,r y��q�����q�a r�T�n�t�����	t�KNOW_M�  |uGvz�SV7 ��z�rs &����>/�/PG/�a��y�MM���{� ���	^r�` (l+/�/',~�$@X�	����@���%�"�4�.0pz�MRM��|-TU�y�c?u;e�OADBANFW�D~x�STM�1 k1�y�4e� �8��̾�?�?�?(OO -O?OqOcOuO�O�O�O �O�O�O&___\_;_@M_�_q_�_�_�72�<8�!�?�`�<�_�_�N�3�_�_
oo�74 9oKo]ooo�75�o�o�o�o�76�o�o��772DVh�78`�����7MA�0���swwOVL/D  �{�/a��2PARNUM � �;]�o��3SC-H*� 8�
����8ω�3�UPD��[��ܵ+�wu_CMP_0r -��0�'�5C��ER_CHKQ�����1�"e�N�`�RqS>0�?G�_MO�?�_��#u_RES+_G�0��{
Ϳ @�3�d�W���{����� ���կ���*�����P��O��8` l�������`��ʿϿ ��`�	���1p)� H�M���phχό����p�������V 1���5�1�!@`y��ŒTHR_IN�R>0/�Z"�5d:�M�ASSG� Z[�M�NF�y�MON_QUEUE ��5��6Ӑ~#tNH�U⌑N�ֲ���END8�����EXE������BE������OP�TIO������PR�OGRAM %���%��߰���T�ASK_I,�>�O?CFG άߞ������DATAu#�&����Ӑ2�%B� T�f�x���5������� ������,>P��INFOu#� �� ������� '9K]o�� ������/lx� � ;���ȀK_�����S&�ENB-�b-&q�&2��/�(G��2�b+� X,		��=�����/��@��P4$�0��99)��N'_EDIT ����W?i?��WER�FL�-ӱ3RGA�DJ �F:A�  �5?Ӑ�5Nј6���]!֐��?�  Bz�W"Ӑ<1Ӑn&%�%O0�8;��50!2��7�k	H��l0�,�{BP�0�@�0��M*�@/�B **:�B�O�F�O2�	�D��A�ЎO�@O�	_,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_�_ o�_o�_�_
o�o.o �ojodovo�o�o�o�o �o�o\XB<N �r����4�� 0���&���J����� ������������ x�"�t�^�X�j�䟎� ��ʟğ֟P���L�6� 0�B���f��������� (�ү$������>� ��z�t��� Ϫ���� ��l��h�R�L�^�DX	���ώ0�� ���t$ :�L��o��
ߓߥ��7PREF� ��:�0�0
~�5IORITYX��M6��1MPDSP0V�:n" �UT��C��6ODUCT��eF:��NFOG[@�_TG�0��J:?�HIBIT_DO�8���TOENT 1��F; (!AF_INE*�����?!tcp����!ud��8�!icm'��N?�kXY�3�F<��1�)� �A�����0�����������'  ]D�h�� ����*>��3���9n"OTf�3>S���2�B�G/�LHC��4�;LFJAB?,  ���F!@//%/7/�5�F��Z�w/�/�/�/�3�&ENHANCE� �2FBAH+d �?�%;����������1�1PORT_WNUM+��0����1_CARTR�E�@��q�SKS�TA*��SLGS6������C��Unothin�g?�?OO�۶0T?EMP �N�"O��E�0_a_seiban|߅OxߕO �O�O�O�O_�O'__ K_6_H_�_l_�_�_�_ �_�_�_�_#ooGo2o koVo�ozo�o�o�o�o �o�o1U@e �v����������Q�<�u�.IVOERSI	�L���� disab�le�.GSAVE� �N�	26�70H771|�h��!�/��9�:�C 	^�4�ϐ����e��͟ߟ���A��9�D�C-Å_y�W 1�������ő����Ǻ�UR�GE� B��r�WAFϠ��-��9�W�����l:WRUP_�DELAY ���=n�WR_HOT %��7��/p���R_NORMAL�O�V�_�����SEM�I��������QSKKIPo��97��xf� =�b�a�sυ�H��ʹ� �ø��������&�� J�\�n�4�Fߤߒ��� ���߲���� �F�X� j�0��|������� �����0�B�T��x��f���������ãRB�TIF�5���CV�TMOU�7�5]���DCRo���� �T�+����B���C�jP>�4J^�9�L�&H͵����jW�ſE����VϦ��<
6�b<߈;܍��>u.�>*��<��ǪP0���2DVh z��������,GRDIO_TYPE  v��/�ED� T_CFGg ��-�BH]��EP)�2��+ ��B�u �/�* ��/�?�/%?=�/ V?�}?�Ϟ?���?�? �?�?�?O
O@O*Gl? qO��8O�O�O�O�O�O �O�O�O_<_^Oc_�O �__�_�_�_�_�_o �_&oH_Mol_o�oo �o�o�o�o�o�o�o" DoIho*j�� �����.3�E� �f� ���x������� �ҏ�*�/�N��b� P���t�����Ο��ޟ��:�+���R'INT� 2�R��!�1G;� i�{��"���8f�0 ��ӫ� �����M�;�q� W�������˿���տ �%��I�7�m��e� �ϑ��ϵ�������!� �E�3�i�{�aߟߍ� �߱���������A����EFPOS1 �1�!)  x���n#������� ������/��S��� w����6�����l��� ����=O����6 ���V�z�  9�]��� �Rd���#/� G/�k//h/�/</�/ `/�/�/??�/�/? g?R?�?&?�?J?�?n? �?	O�?-O�?QO�?uO �O"O4OnO�O�O�O�O _�O;_�O8_q__�_ 0_�_T_�_�_�_�_�_ 7o"o[o�_oo�o>o �o�oto�o�o!�oE W�o>���^ �����A��e�  ���$�����Z�l��� ��+�ƏO��s�� p���D�͟h�񟌟� '�ԟ�o�Z���.� ��R�ۯv�د���5� ЯY���}���*�<�v� ׿¿����Ϻ�C�޿�@�y��e�2 1� q��-�g�����	�� -���Q���N߇�"߫� F���j��ߎߠ߲��� M�8�q���0��T� ��������7���[� ����T�������t� ����!��W��{ �:�^p�� A�e �$ ��Z�~/�+/ ���$/�/p/�/D/ �/h/�/�/�/'?�/K? �/o?
?�?.?@?R?�? �?�?O�?5O�?YO�? VO�O*O�ONO�OrO�O �O�O�O�OU_@_y__ �_8_�_\_�_�_�_o �_?o�_co�_o"o\o �o�o�o|o�o)�o &_�o��B� fx��%��I�� m����,���Ǐb�� �����3�Ώ���,� ��x���L�՟p����� ��/�ʟS��w����<�ϓ�3 1��H� Z������6�<�Z��� ~��{���O�ؿs��� �� ϻ�Ϳ߿�z�e� ��9���]��ρ���� ��@���d��ψ�#�5� G߁�������*��� N���K����C��� g��������J�5� n�	���-���Q����� ����4��X�� Q���q�� �T�x� 7�[m�// >/�b/��/!/�/�/ W/�/{/?�/(?�/�/ �/!?�?m?�?A?�?e? �?�?�?$O�?HO�?lO O�O+O=OOO�O�O�O _�O2_�OV_�OS_�_ '_�_K_�_o_�_�_�_ �_�_Ro=ovoo�o5o �oYo�o�o�o�o< �o`�oY�� �y��&��#�\� ������?�ȏ����4 1�˯u����� ?�*�c�i���"���F� ���|����)�ğM� ����F�����˯f� ﯊�����I��m� ���,���P�b�t��� ���3�οW��{�� xϱ�L���p��ϔ�� �������w�bߛ�6� ��Z���~�����=� ��a��߅� �2�D�~� �������'���K��� H������@���d��� ��������G2k �*�N��� �1�U�N ���n��/� /Q/�u//�/4/�/ X/j/|/�/??;?�/ _?�/�??�?�?T?�? x?O�?%O�?�?�?O OjO�O>O�ObO�O�O �O!_�OE_�Oi__�_ (_:_L_�_�_�_o�_ /o�_So�_Po�o$o�o�Ho�olo�oۏ�5 1����o�o�olW ��o�O�s�� �2��V��z��'� 9�s�ԏ��������� @�ۏ=�v����5��� Y��}�����۟<�'� `��������C���ޯ y����&���J���� 	�C�����ȿc�쿇� ϫ��F��j�ώ� )ϲ�M�_�qϫ���� 0���T���x��u߮� I���m��ߑ����� ���t�_��3��W� ��{������:���^� ����/�A�{�����  ��$��H��E~ �=�a��� ��D/h�' �K���
/�./ �R/��/K/�/�/ �/k/�/�/?�/?N? �/r??�?1?�?U?g? y?�?O�?8O�?\O�? �OO}O�OQO�OuO�O�O"_t6 1� %�O�O_�_�_�_�O �_|_o�_o;o�__o �_�oo�oBoTofo�o �o%�oI�om j�>�b��� ����i�T���(� ��L�Տp�ҏ���/� ʏS��w��$�6�p� џ���������=�؟ :�s����2���V�߯ z�����د9�$�]��� �����@���ۿv��� ��#Ͼ�G�����@� �ό���`��τ�ߨ� 
�C���g�ߋ�&߯� J�\�nߨ�	���-��� Q���u��r��F��� j������������ q�\���0���T���x� ����7��[�� ,>x���� !�E�B{� :�^����� A/,/e/ /�/$/�/H/ �/�/~/?�/+?�/O?<5_GT7 1�R_�/ ?H?�?�?�?�/O�? 2O�?/OhOO�O'O�O KO�OoO�O�O�O.__ R_�Ov__�_5_�_�_ k_�_�_o�_<o�_�_ �_5o�o�o�oUo�oyo �o�o8�o\�o� �?Qc��� "��F��j��g��� ;�ď_�菃������ ˏ�f�Q���%���I� ҟm�ϟ���,�ǟP� �t��!�3�m�ί�� 򯍯���:�կ7�p� ���/���S�ܿw��� ��տ6�!�Z���~�� ��=ϟ���s��ϗ� � ��D������=ߞ߉� ��]��߁�
���@� ��d��߈�#��G�Y� k�����*���N��� r��o���C���g��� ��������nY �-�Q�u� �4�X�|b?t48 1�?);u ��/;/�_/� \/�/0/�/T/�/x/? �/�/�/�/[?F??? �?>?�?b?�?�?�?!O �?EO�?iOOO(ObO �O�O�O�O_�O/_�O ,_e_ _�_$_�_H_�_ l_~_�_�_+ooOo�_ soo�o2o�o�oho�o �o�o9�o�o�o2 �~�R�v�� �5��Y��}���� <�N�`��������� C�ޏg��d���8��� \�埀�	�����ȟ� c�N���"���F�ϯj� ̯���)�įM��q� ��0�j�˿��ￊ� Ϯ�7�ҿ4�m�ϑ� ,ϵ�P���tφϘ��� 3��W���{�ߟ�:� ����p��ߔ���A� ���� �:����Z� ��~�����=���a����� �����MA_SK 1����������XNO � ���� MOT�E  �R_C�FG �Y�����PL_RANG�UP���OWE/R ��� ��A��*SYST�EM*P�V9.3�044 �1/9�/2020 A� � ���RE�START_T �  , $F�LAG� $DS�B_SIGNAL�� $UP_C�ND4���R�S232r �� $COMM�ENT $�DEVICEUS�E4PEEC$P�ARITY4OP�BITS4FLOWCONTRO3?TIMEOUe6�CU�M4AUX�T��5INTER�FACsTATU��HCH� t $OL�D_yC_SW �'FREEFR�OMSIZ �A�RGET_DIR� 	$UPD�T_MAP"� T�SK_ENB"E�XP:*#!jFA�UL EV!�R�V_DATA�_  $n E��   	$VAL�U�! 	j&GR�P_   �{!A  2 ��SCR	�� �$ITP_��" $NUMΞ OUP� �#TO�T_AX��#DS}P�&JOGLI�FINE_PCdn�OND�%$�UM�K5 _MIiR1!4PP TN?8�APL"G0_EX�b0<$�!� 814�!P=Gw6BRKH�;&{NC� IS �  �2TYP� �2�"�P+ Ds�#;0BS�OC�&R N�5DU�MMY164�"S�V_CODE_O�P�SFSPD_�OVRD�2^L�DB3ORGTP; LEFF�0<G� �OV5SFTJRUNWC!SFpF5%3oUFRA�JTO��LCHDLY7R�ECOVD'� WaS* �0�E0RO���10_p@  � @��S NVE�RT"OFS�@C� "FWD8A�D4A��1ENABZ6�0T�R3$1_`1FD}O[6MB_CM�!zFPB� BL_M��(!2hRnQ2xCV�"�' } �#PBGiW|8A�Mz3\P��U�B�__�M�P�M� �1�AT�$CA� �PD�2��PHBK+!:&aI�O�4 eIDX+bPPAj?a$iOd�7e�U7a�CDVC_DBG"�a;!&�`��B5�e1�j�S�e3��f�@ATIO� ���AU�c� �S�AB
0Y.#0�D���X!� _�:&S�UBCPU%0S�IN_RS�T, 1�N|�S�T!�1$HW_C1�"]q.`�v��Q$AT! � �_$UNIT�4�p>�pATTRI= �r�0CYCL3NE�CA�bL3FLTR_2_FI9a7�c�,!LP;CHK�_�SCT>3F_ƥwF_�|8��zFS8+�R�rCHAGp�py��R�x�RSD�@`'�1E#&7`_T�X�PRO�`@S�EMOPER_0�3Tf��]p� f��P�DI�AG;%RAILAiC�c4rM� LO�04�A�65�"PS�"�2� -`�e�SPR�`S&.  �W�Ctaf�	�CFUNC�2~�RINS_T.!`(�w��� S_� ��0�P�� 	d��W�ARL0bCBLCUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!��8�3�TID�S��!�� $CE_RIYA !5AFDpPC�~��@��T2 �C�9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@HRgDYOL1	PRG8��H��>1(�ҥMUGLSE =#Sw3��$JJJ6BKGFK�FAN_ALML�V3R�WRNY�HGARD�0+&_P "B��2Q���!�5_�@�:&AU�Rk��TO_SBRvb��� �ƺ�pvc�޳MPINF�@�q�)���'REG'd~0V) 0R<�C�1DAL_ \2sFL�u�2$MԐ (�#S��P� `�gśCMt`NF�qsO�NIP�qEIPPs 9a$Y���! �"�!7� �o3EGP��#�@��AR� �c�52p�����|5AXE�'wROB�*RED�&�WR�@�1_=��3S�Y�0ѥ0_�Si�WcRI�@�ƅpST@�#��0*@� �q	���3��� B� �A��3�]D�POTO�� �@ARY�#��!��d̒!1FI�0�$�LINK��GTH��B T_���Ar��6�"/�XYZ+":9�7G�OFF�@�).�"���B� l�����A3$ ��FI@�p���4�4l��$_Jd�"(B�,a������8�"q�����2�Ck6DUR��]94�TURT�XZ��N����Xx��P��FL/�@s��l�P���30�"Q 1J� K
0M:$�53]q�7�SuD�Sw#ORQ�Ɇ�!�����Q7��0O[�ND�=#�!#�1'OVE8��M� ��R��R��Q!P0.!P! OAN}q	� R����990� �br J9V����v�!SER1��	8�E�@Hn D�A��p�����Ă���v�AX �C�"��`�q�s� ��0~3�~F��~e�~�~E�~1 ��~Ҡ{Ҡ�Ҡ� Ҡ�Ҡ�Ҡ�Ҡ��Ҡ�Ҡ�!)DEBU}s$x�����!R*�AB�a8Ar2V`|r 
�" �c���%�Q7�7�1 73�7F�7e�7�7E�������L�AB����yp�cG�RO�p��}��PB_ҁ ��̓��ð�6��1���5���6AND ��8p�a3���-G �Q����AH�PH�p�2�NTd��Cs@VE�L؁�}A��F�S�ERVEs@�� i$����A!�!�@POR}�KP�иA����@���	  �$�BTRQ�
��CH��@
�G��2	��Eb��_  qlb��Q�ERR��RI�P�@�FQTO	Q�� L�}��YV
ĀG�E%�\���A�RE�  ,h�A�EP
�RA�Q? 2 d�R7cs��T�@ ��$F ׂ��m���B�OC��P  }8[COUNT����@�SFZN_wCFG�A 4�p%��rT\zs�a�#`p�Jp b ��(a�� �� MGp+����`0�OGp�eFAq����cX8еk�ioQ�¤'ѴDp8�Pz���SHELA�-b� 5��B_wBAS\RSR$Ɗ`�2�S��L�!p1T�W!p2Dz3Dz4DzU5Dz6Dz7Dz8�WqROO���P�1�3NL�� �AB�C
�n"pACK�&IN�P	T+�W�U��	�k��y�_PU8�~�|�OU�CP��%�s�Vl����YTPFWD_KcARKQ-�:PRE�D��P����QUE�$�Ā9 )���~���I U��#s/���@�/�SEM1ǆ1�An�aSTY�tSO����DI�q��Qc��X_TM9�MANsRQ �/�END���$KEYSWI�TCH2�G����H}E)�BEATMz�PE��LEJR���0Jx�UF�F��G�S��DO_HOM��Olz��pEFPR��PSbJі��uC��O��<7P�QOV_M��}�c�IOCM���1�.� uHK�� �D,�&�a`U2R��M���a�r +�FORC�*�WAR��� uOM��  Q@�$�㰰U��P�Q1��g���3��4�1T�B�POW�Lz��R�%�UNLO�0T��ED��  ��SNP��S.b �0N�ADDa`z��$SIZ*�$V�A�0�UMULTI�P�r���Az�? � $��Hƒ���SQc�1CFP�v�FRIFr�PS�w���ʔf�NF#�ODBUx�R@w������F��:�IAh�����������S"p�� g�  �cRTE��\�SGL.�T�x�&C`Gõ3a�/�S'TMT��`�P�����BW9 0�SHOW�h�qBANt�TP o���E������PmV_Gsb ��$PC�0�PoF�Bv�P��SP��A��p���`VD��rb�� �+QA002D.ҝ�6ק�6ױ��6׻�6�54�64�7�4�84�94�A4�B�4و�6ׇ17�}�6�F 4� ��@�����Z��T��t�1��1��1��U1��1��1��1��U1��1��1��23�U2@�2M�2Z�2g�U2t�2��2��2��U2��2��2��2��U2��2��2��33٨���M�3Z�3g�3�t�3��3��3��3���3��3��3��3���3��3��43�4�@�4M�4Z�4g�4�t�4��4��4��4���4��4��4��4���4��4��53�5�@�5M�5Z�5g�5�t�5��5��5��5���5��5��5��5���5��5��63�6�@�6M�6Z�6g�6�t�6��6��6��6���6��6��6��6���6��6��73�7�@�7M�7Z�7g�7�t�7��7��7��7���7��7��7��7���7��7���VPzv�U�B �@��09r
�@V���A/ x �0R���+  �BM�@RP�`�4Q_�PR�@[U�A�R��DSMC��E�2F_U��=A��YS�L�P�@ �   �ֲ>g�������<iD��VALU>e�p�L�A�HFZAID_YL���EHI�JIh�?$FILE_ ��D��d$ǓB�XCSA��Q h�0!PE_BLCKz�.RI�>7XD_CPUGY!�@GY�Ic�O
T�`Y.���R  � �PW`�p���QLAn�S�Q�S�Q�TRUN_FLG�U �T�Q�TJ��U�Q�T�Q��UH��T`�T�T�2L�_LIz� w �pG_O}T�P_EDIU�c��/`�`7c ?b�ة�pBQh����T�BC2 �! ��%�>��P��a�7aFT�τ�d݃TDC�PA�N`�`M�0�f�a�gTH��U��d�3�g�R�q�9�ERVE Ѓt݃t	��a�p��` "X -$EqLENЃRt݃�Ep�pRAv��Y@WI_AtS1Eq�D2�w�MO?Q�S���pI��.B�A�y�4Ep�{DyE�u��LACE ��CCC�.B��_M�A��v��w�TCV�:��wT,�;�Z��P���s�~��s�JJ�A�M����J����uā�uQq2�ѐ���݁�s�JK��VK������	�b��J����JJ�;JJ�AAL�<� �<�6��:�5�cm��N1a�m�,��DL²p_\�Ű�1ApCF�
�# `�0GRO�U�@J�Բ��N�`C�^�ȐREQUIRrÀEBUu�Aq��7$T�p2"��Bpp薋a	��d$ \?@�qhAPPR��CL�B
$H`N;�CL	O}`K�S�e`��u��.I�% �3�M�`�8l��_MG񱥠�C �"P����&���B{RK��NOLD����RTMO6a�ޭ��J6`�P>��p���p��pZ��pc��p6+�7+�<��QAq�d&� �lr���������PATH ��������qx�����9%0A��SCAub��l<���INDrUC�p��q�C�UM�Y�psP����A q/��/�E�/�PAYL�OA�J2L�0R'_AN�ap�L�Pz��v�jɆ���R_F2�LSHRt��LO�{�R�������ACRL_�q�����b�rd�H�@B$H��^"�FLEX>�.`;BJ�f' P(��o��o+�p�aJDu( :Qcv�p�׀��fe��po��|F1���-������]�E��*�<� N�`�r�����4�Q��� ����A�c���ɏۏ���T��2�X:A��� ���������)� ;�?�H�6�Z�c�u���t��?qJ��) ��``��˟ݟ�`�0ATF�𑢀EL���a���J�(��JE۠C3TR��A�TN�1��HAND_VB�B>ѯ@�* $���F2���d�CS�WR����+� $$M�����0ˡ�@ڡ������A�@ g����A)��A���@
˪A٫A� ��`P�˪D٫D�PȰG�P�)STͧ�!ک�!N�DY�P9���� #%��Fp���Ѫ���i� ���������P3�<��E�N�W�`�i�r�  ���, ��ԓ�� n�5m��1AS�YMص.@�ض+A������_`��	� ��D�&�8�J�\�n�Ju�&��ʧC�I��.S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R�� &T��3TWV�͢���&���ߪU��/�7� ̢1�`HR`ta-0��QQ�1�DI���O�T��P��. ; *"IAA*���$a`G�2C2cJ��`_�H���P / � �ME�� Mb�R4AT�PPT�@� ��ua���P�l@zh�a�iT�@�� $�DUMMY1E�o$PS_D�RF���P$�f3�FL�A��YP���b}c?$GLB_T��U�uu`1��0��EQa0c X(���ST�����SBR�PM2�1_V��T$SV_ER��O_@KscsSCLpKrA��O'b��PGL�@EW��1s 4��a$Y|�Z|W�s怯��A\N`� ��sU�u�2 ��N�p�@w$GIU}$�q 1�s�p���3 L���v^B}$�F^BE�vNEARʖ�NK�F8���TAsNCK��QJOG���� 4��$JOINT�� x��q�MSET��5  ��wE�H�� S�@��� ��6�  �MU��?���LOCK_FO����PoBGLVHGL�TEST_XM>�N��EMPt�[��r̀$U�Гr��#22���s,�3���4Ҁ,�1MqCE���s�M� $KAR��M>�STPDRA�pj��a�VEC��{�e�I�U,�41�HEԀT�OOL㠓V�R�E��IS3����6�N�A�ACH���5���O�}c�d3����pSI.�  @�$RAIL_BO�XE��ppROB�O��?�pqHOW�WAR*���`�ROLM�bB���S�p�
�5���O_F� �!ppHTML5�Q�����0�r�ڑ��7m���R
��O��8m��v�z��ЍtOU��9 tpp(�14A�̀���PO֡%PIP��N��
�ڑS�,������CORDED0Ҁް̠5�XT��q�)HbP� O4` �: D pOB P!"Ҁ{�j��cpj��^@$SYSj�ADqRFa�Pu`TCH�� ; ,��ENT�RZ�Aف_�t״x���QVWVAPa?< � p��r��UPREV_RT~]1$EDIT�_VSHWR�7v(;���q�@D_`#�R�+$HEA�DoA�Pl�A$�K�E�q�`CPSPD.��JMP��L�U� R��d=r�O�϶�I�S#CiNEx��$_TICK�ʅAMX�~���HN-q> @t�������_GP��[�S3TYѲ�LOq�����Ҩ�?�
�G�ݵ%$���t=7pS !$Q��da�e�!`�fP�0�SQU�d� ��b�ATERC�y`|�pS�@ �pCp����d�b%Oz`mcO�IZ�d4�q�e�aPRM��a�8����PUQH�_�DO=�ְXS��KN�VAXIg�f�1�UR� ��$#�Е�d�� _����ET��QPۂ���5f�F�7�g�A�!�1�d9��2;���R|Al�о�� �#��5��#��#� )#�)i�>'i�N'i� ^&{����){����2��	C����C��WOiO{O��D��TSSCp oB hppDS(��k��`SP`�AT�L �I���¼bA_DDRES��B'��SHIF��"�_2+CHF`��I&p���TU&pI� }Cm�CUSTO��*	aV��IbDȲ�,��0
�
��V8�X�R`E \����A�f�7��tC�#�	���F��irt�T�XSCREEl�Fz�P��TINA�s�p��t�q���0G T��fp,⧱eq�Bp&uᦲu�$#�RRO'0R�F`}�!Cdv �UE��H ��0����`S�q��RSM�k�UV����V~!�PS_�s�&C�!�)�'�C��Cǂz"� [2G�UE�4Ib�vr�&8�GMTjPL�DQ��Rp�z�BB�L_�W�`R`J ��f�>2O�qJ2L�E�U3"�T4RI;GH^3BRDxt�OCKGR�`�5TW�|�7�1WIDTH��H�Bb�a�a��	��UIu�EY��QaK� d�p��A�J�
�4�BACKH��b�5�|qX`FOD�GL[ABS�?(X`I�˂$UR(�9@����0^`H4! L 	8�QR�_k��\B_`R�p͂����a�IA)O�R`M��w0�Uj0�CRۂM�LUqM�C��� ERV��	`�0P<��4NV`��GE=B#���]�t��LP�E��E��Z)�Wj'Xz'XԐ&Y5*$[6$[7$[8	R��@�3�<���fԑŁ�S��M�1USR��tO <��^`U��r�rFO
�rP�RI��m����PT�RIP�m�U�NDO��P�p ��`m�4���#����� QWB�P7�G �s�Tf�H�RbO	S�agfR��:">c��.qR��s�~�b*�~�#�UQ.qS�o�o�#8R)�>cOFF���p�T� �cOp �1Rppt/tSppGU��P.qx�JsETwn�1SUB*� f�_E_EXE��V��v>cWO>� U�`^g��WA'��P�q�!@� V_DB8�s�p�BSRT�`
�aV�Q�r��OR�N�uRAU��tT��ͷ�q_���W |�%�͸OWNA`޴�$SRCE � ��Dx��\��MPFIA�`��ESPD��� ���C���Gƒ�)�5���!X `�`�r޴���COP�a$��C`_w�������rCT�3�q���qƒpp��@� Y"?SHADOW�ઓ~@�_UNSCA��8@��4M�DGDߑ��OEGAC�,Me��G�Z (0N�O�@�D<�PE�B&��VW씪�G���!�[ � ��VE8E#��ڒANG�$���c薴cڒLIM_X�c��c� �����#��`� 퐾�VF<� �s�VCCjв�5\ՒC{�RAlצ����RpNFA���%�E��Z`G̭ ^0[�C`DE8Ē��� STEQ1�� �@�ꁻ@I��`+0����`����P_A�6�r���K��!]G� 1Ҡ������\��сCPC�@]�D#RIܐ\�͑V#Ѐ����D�TMY_UBY�T���c��F!����Y��$���P_hV�y��LN�BMQ1�$��DEY��E�X�e��MU��X�M� US�!���P�_R����P� ߖG��PACIr�ʐf� ᔟ��c�´c���#�!EqB��a.2B���N�^ ܀Gΐ!P���40C�R~``�A_�0�@3!�1zr	�e�R�SW��p�00H��S�6�O�Q�1A� 4X�#�E�UE��00Y)�D�HKJ�`�@�p���U� �EAN�ٖp�pXՆ`C��MRCV�!a ���@O��M�pC�	p��s����REF*7 
��������/��P�ڀ@���@��b��֗�_ Y��ژ��ۣ��Q$3�������AC��$b �����%���Q��$GROU� �c������ʠ]��I2^`0��U` 0_��I,�o � ULա`2��C&�rAaB�?�NT����$����A���Q��K�L����õ���A���Q��T a$c� t�`MD�p8�H�U���SA��CMPE F  _�Rr�p@����9XS	��VGF/�b#_d, &�@M�P^0۰UF_C !���z �ROh0"+��p�@���0C�UREB����RI��
IN �p�����d��d�,�ca�INE�H�y��0V�a-�걗�3�W�������C��i�LO�}�z�@0�!�QNSI��݁����c$&�c$&.�X_PuE-YW+Z_M�ڒW�I�$�" �+�R�'rRSLre� �/�M
`�RE�C7�Gd�۰�� �ҭ�q����u��� �������S_P�V�nP ��IA�vf� �~pHDR�p�pJO�P��_$Z_UP��a_LOW�5�1J�dA���LINubEP�?�tc_i�1�1���@��G1@��V�xg{ 5X�PATHP= X�CACH$��]E��yI�A��{�C�)�ID3FA�ETD��H��$HO�pO�b@�{�d6�F����<��p�PAGE�䁀�VP�°�(R_SI	Z��2TZ3�-X�0U̲q�MPRZ��IM5G���AD�Y��MRE��R7WGP���8�p��ASYN�BUF�VRTD��U�T7Q�LE_2�D-��U��`CҡU�1��Qu��UECCU��VEM��]EDb�GVIRC�Q�U�S��B�Q�LA��p�N�FOUN_�DIAuG�YRE�XYZ�cE�WѴh8�dpq2a`T��2�IM�a�V�|be��EGRABBr��Y�a�LERj��C4���FC-A�65a04x��7u$� BE���h��`�CKL�AS_@l�BA��N@i�  G��T��� @�ݲմ$BAƠwj A�!q�eb��uTYS p�H����2��I�t:bt�f��B)�EVE�����PK���fx��G�I�pNO��2����rHO����k � ���
8�Pi��S�0ޗ��RO��AOCCEL?0=���VR_�U7@�`��2�lp��AR��PA���̎K�D��REM_�But � #�JM�X �l�t�$S�SC�U�ҫ2�OG��QN@m � �S�P�NS���LEX�vn T�ENA�B 2�W@��FLDRߨFI�P�t�ߨ�(Ğ�1��P2>HFo� ���V
Q MV_PI ��8T@󐉰�	F@�Z�+�#��`8�8#��GAB�Ε�LOO��JCqBx��w"SCON(P�PLANۀ�Dp��3F�d�v�9PէM ��Q ;����SM0E� ɥ�8ɥWb72$`d<�8T��,`RKh"�ǁVANC��FR��VR_Ou N@p (�-#<#c��c�2
�R_A/�N@q 4������`	�^�8�0w�N@r hn��8�1^�&OFF`|�ap�`��`�DEA�Y
�P,`SK�DMP6�VIE��2q �w��@���rs < !{���4���r{7���D���}qCU�ST�U��t �$G�TIT1�$PR\��OPT<ap ��VSF�йs�u�p�0`r&�.M�SMOwvI�|��ĄJ�����eQ_$WB��wI���� @�O3�@�XVRx�xmr��T����ZABC��y �op����)�
e�Z�D$�CSCH��z Lu����`�2�%P0C ��7PGN ��x<��A��_FUNH���@ˑZIPw{,I��LV,SL��~��� �ZMPCF���|��E����X�DMY_LNH�=�C��� ��} $x�A� ]�CMCM� EC,SC&!��P��? $J���DQ������������±�_�Q,2����UX|�a\�UXEUL� �a������(�:�(�<J���FTFL��w�C��~Zp+�6�S ﰑ�Y@Dp�  8 $�R�PU��> EIGH����?(�iֱ�qb���et� �a�����$B�0�0@�}	�_SHIFD3�-�RVV`Fcв�		$5��C�0��&!������b
�sx�uMD�TR��V̱����SPH���!�� ,�������	��4A�RYP��%������%�A�"��%!  �H�(UN0���"�2X����� �q0GSPDak����P��O��`��0�āЯ�}"!NGVER`q7 iw+�I_AIRPUR�GE  i C i/�F`E�Tb�; �+  � h2ISOLC  �,E�"�!A��!�%d��P+�_/*OB���Dm�?@�!�H771  34n?�?�9� `�E�/#�)x� S232Γ� 1i� �LTEk@ PENDA�341 1�D3<*? �Mainte�nance CoKns B�? F"O�,DNo Use MJOOnO�O�O�O�O2�2NPO;/" 159%�1CH=����-Q		9Q_!�UD1:___RSMAVAIL/��/%�A!SR  �+��H�_�P1�oTVAL.&����P(.�YVL�}� 2�i�� D��P��/`oVPNo�o rci�o�g�o�o�o�o �o*,>tb �������� �:�(�^�L���p��� ����܏ʏ ��$�� H�6�X�~�l�����Ɵ ���؟�����D�2� h�V���z�������� ԯ
���.��R�@�b� d�v�����п����⿀��(�N�<�r�i��$SAF_DO_PULS. jQp�����CA� �/%��&0SCR ��`X��A�A�
	14�1IAIE��@� S�wo%�7�I�[� m��ߣߵ������߬���GS��2H%��0�d%�@�rb��� @�"k�}��T�h� J`����_ @��T�7 �����#�0�T D��0�Y�k�}� �������������� 1CUgy�O�Ef�����  �5;��o�� 1p�U�
�t��Di��������
  � ��*������gy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�?��?�?OO%O7O<A� ��`OrO�O�O�O�O�O �O�O?O�_._@_R_ d_v_�_�_�_�_�Q _�R0MJTo!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏJO ��'�9�K�]�o��� ����_ɟ۟���� #�5�G�Y��_�U�_�� ������ϯ���� )�;�M�_�m������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T�f�;�?�q߮��� ��������,�>�P� b�t�������������������Y��	12�3456781�h!B!����F������� ����������  ��;M_q��� ����%7 I[l*���� ���//1/C/U/ g/y/�/�/�/n��/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O �/)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_O_�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�op_�o �o�o/ASe w������� ��o+�=�O�a�s��� ������͏ߏ��� '�9�K�]�������� ��ɟ۟����#�5� G�Y�k�}���������s�կ�w����0�L�CH  B}pw�   �=��2�� }� =�
���  	�o�ί��ǿHٿ���r������ @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖ�%Ϻ����� ����&�8�J�\�n� ��������������"�Q�*�����;��<M���D���  �]�w�*�Z�|����t  d�����*�`*��$S�CR_GRP 1�*P3� �� �*�� 6�	 _�
 ��<�+*�'U8C|@��y�yD� W�!�y��	M-10i�A/7L 1234567890���� 8��MT� � �
�	L��Y	Č� N
����Y���y�
M_	P������ ,��H�
 ���1/@@A/g/y/H�ߙ!T/��/P/�/3��+���/B�S��,?*2C4&9Ad�R?  @s�j5N?�7?��7&2R��?�}:&F@ F�`�2�?�/�?�?OO -OSO>OwObO�O=j1��2�O�O�O�O�DB� �O�O;_&___J_�_n_ �_�_�_�_�_o�_%o��5j�eSgxo6����uo�o�b�1j17��.�oh0�4j9j9B� w�$Y̯@HtA�Nhcu�/�%Ipp�drsq ����z�q�x� �.� (&�*�2� D�V�oz�e��������ECLVL  Ψ���iqpQ@���L_DEFAU�LT ���s�փHOT�STR⍝q��MI�POWERF���H���WFDO�� �RVENT 1ɁɁ�� L!DUM�_EIP�����j�!AF_INEx‧���!FT}��֞����!-/� ���F�!RP?C_MAING�)�q�5���Y�VISb��t����ޯ!TP&ѠPUկ��dͯ*��!
PMON_POROXY+���e��v��D���fe�¿!�RDM_SRV�ÿ��g���!R�,*ϑ�h��Z�!
�[�M����iIϦ�!RLSYNC�����8����!R3OS|���4��>��!
CE�MTC�OM?ߓ�k-ߊ�!=	S�CONS�ߒ��ly���!S�WA'SRCݿ��m��"�;!S�USB#�n�n�!STMC��o]����� ѳ����,���P�V��ICE_KL ?�%d� (%S?VCPRG1S���"��2������3����"��4������5"��6;@��7ch������9�� ��%�������� 0����X����� -���U���}� �� /���H/��� p/���/��F�/�� n�/��?��8? ���`?��/�?��6/ �?��^/�?��/X�j� ��q���#OhO��lO�O {O�O�O�O�O�O�O _ 2__V_A_z_e_�_�_ �_�_�_�_�_oo@o +odoOo�o�o�o�o�o �o�o�o*<` K�o����� ��&��J�5�n�Y����}���ȏ���^�_�DEV d���MC:�4����GRP 2�d�
@�bx 	� 
 ,V��o�u�[������ �����ٟ���:�L� 3�p�W�������ʯ�� � �W�$�ۯH�Z�A� ~�e�������ؿ���� ���2��V�=�zό� sϰ�����ϝ�
��� .�@�'�d�K߈ߚ߁� �ߥ����������<� #�5�r��ϖ����� ��������&��J�1� n���g����������� ����"4��X| �u����� �0)fM�q ����;�/� >/%/b/t/[/�//�/ �/�/�/�/?(??L? 3?p?W?i?�?��?�? �? O�?$OOOZOAO ~OeO�O�O�O�O�O�O _�O2__V_h_�?�_ C_�_�_�_�_�_
oo o@o'odoKo]o�o�o �o�o�o�o�oo_ NrY���� ����&��J�\� C���g�������ڏ�d ��	ȏ����5� �Y�D�}���%�x���������ʑ v�ʕڟ�ҟ���,� �P�^�����ƙF��� ��ԯ¯����.�p� U������v�����п ���6�\�-�l��`� Nτ�rϨϖ������ 2ϼ�&߸�6�\�J߀� nߤ�����
ߔ����� "��2�X�F�|�ߣ� ��l����������� .�T���{���D����� ��������\�AS 
,t���� �4X�L:\ ^p����0 �$//H/6/X/Z/l/ �/��//�/�/�/ ? ?D?2?T?�/�/�?�/ z?�?�?�?�?O
O@O �?gO�?0O�O,O�O�O �O�O�O_ZO?_~O_ r_`_�_�_�_�_�_�_ 2_oV_�_Jo8ono\o �o�o�o�o
o�o.o�o "F4jX��o ��~�z��� B�0�f�����V��� ��Џҏ���>��� e���.���������̟ Ο���X�=�|��p� ^���������ȯ�D� �T��H�6�l�Z��� ~�����ۿ���Ϡ� �D�2�h�Vό�ο�� �|�����
����@� .�dߦϋ���T߾߬� ��������<�~�c� ��,��������� �D�)�;������\� �����������@� ��4"DFX�| ������0 @BT���� z��/�,//</ ���/�b/�/�/�/ �/?�/(?j/O?�/? �??�?�?�?�?�? O B?'Of?�?ZOHO~OlO �O�O�O�OO�O>O�O 2_ _V_D_z_h_�_�_ �O�__�_
o�_.oo Ro@ovo�_�o�ofo�o bo�o�o*N�o u�o>����� ��&�hM����� n���������ȏ��@� %�d��X�F�|�j��� �����,���<�֟0� �T�B�x�f���ޟï ��������,��P� >�t�����گd�ο�� ���(��Lώ�s� ��<Ϧϔ��ϸ����� ��$�f�Kߊ��~�l� �ߐ��ߴ���,��#� ������D�z�h��� �����(���
�,� .�@�v�d������� � ������(*< r�����b��� �$z�q� J������/ R7/v /j/�z/�/ �/�/�/�/*/?N/�/ B?0?f?T?v?�?�?�? ?�?&?�?OO>O,O bOPOrO�O�?�O�?�O �O�O__:_(_^_�O �_�_N_p_J_�_�_�_ o o6ox_]o�_&o�o ~o�o�o�o�o�oPo 5to�ohV�z� ���(�L�@� .�d�R���v����� �$�����<�*�`� N���Ə���t�ޟp� ���8�&�\����� L�����گȯ�� ��4�v�[���$���|� ����ֿĿ��N�3� r���f�Tϊ�xϮϜ� ���������Ͼ�,� b�P߆�tߪ������ �������(�^�L� ���ߩ���r����� � ����$�Z������ J������������� b���Y��2�z� ����:^� R�b�v��� �6�*//N/</ ^/�/r/�/��//�/ ?�/&??J?8?Z?�? �/�?�/p?�?�?�?�? "OOFO�?mOO6OXO 2O�O�O�O�O�O_`O E_�O_x_f_�_�_�_ �_�_�_8_o\_�_Po >otobo�o�o�o�oo �o4o�o(L:p ^��o�o�� � �$��H�6�l���� �\�ƏX�֏��� � �D���k���4����� ��ҟ����^�C� ���v�d��������� ί��6��Z��N�<� r�`����������� ��̿���J�8�n�\� ��Կ������������ ���F�4�j߬ϑ��� Z��߲���������� B��i��2����� ��������J�p�A��� �t�b����������� "�F���:��Jp ^�������  6$FlZ� ������/� 2/ /B/h/��/�X/ �/�/�/�/
?�/.?p/ U?g??@??�?�?�? �?�?OH?-Ol?�?`O NOpOrO�O�O�O�O O _DO�O8_&_\_J_l_ n_�_�_�O�__�_o �_4o"oXoFoho�_�_ �o�_�o�o�o�o0 T�o{�oD�@ �����,�nS� ����t��������� Ώ�F�+�j��^�L� ��p�������ܟ�� B�̟6�$�Z�H�~�l� ���ɯۯ�������� 2� �V�D�z���������$SERV_MAIL  ����ƸOUTP�UTո��@ʴRV 2vj�  � (r�x��<�ʴSAVE����TOP10 2}� d � �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z�`l�~���j�n�YPY��ǳFZN_CFGw j���=��J���GRP �2��g� ,B�   A �D;� B �  �B4=�RB2�1I�HELL��!j�e�)�*����>�%RSR�� ����&J 5G�k�������.�  ���/>/P/"\/ ��X/z"{ �U'&"2�dh,g-�"�EHK 1S �/�/�/�/#?L? G?Y?k?�?�?�?�?�? �?�?�?$OO1OCO??OMM S�O�DFTOV_EN�Bմ�e��"OW_?REG_UI�OȲ�IMIOFWDL�~@�N�BWAIT�B�)��V��F��YTIM�E��G_VA԰_�A_UNIT�C~VeɻLC�@TRY�G�e�ʰMON_ALIAS ?e�I%�he��oo&o 8oFj�_io{o�o�oJo �o�o�o�o�o/A Sew"���� ����+�=��N� s�������T�͏ߏ� ����9�K�]�o��� ,�����ɟ۟ퟘ�� #�5�G��k�}����� ��^�ׯ�����ʯ C�U�g�y���6����� ӿ忐����-�?�Q� ��uχϙϫϽ�h��� ����)���M�_�q� �ߕ�@߹������ߚ� �%�7�I�[���� �����r������!� 3���W�i�{���8��� ����������/A Se����� |�+=�a s��B���� /�'/9/K/]/o// �/�/�/�/�/�/�/? #?5?�/F?k?}?�?�? L?�?�?�?�?O�?1O COUOgOyO$O�O�O�O �O�O�O	__-_?_�O c_u_�_�_�_V_�_�_��_ooc�$SM�ON_DEFPR�OG &����Aa &�*SYSTEM�*obg $J�O0dRECALL� ?}Ai ( �}bo�o�o�o�o�o� })copy� mc:dioc�fgsv.io �md:=>10.�109.3.62:2008	Wi�{{3rfrs:�orderfil�.dat vir�t:\temp\4{6Bp����q+�v*.d��{��Z�l�~�x
xyz�rate 61 �(�:�L�ݏ��u���� ��̏]�o����u6��xmpba�ck��O����� [}-sdb%�*���*�̟]�o���u1x��:\&���8�H�Q�P����p2��a�� ��N�Яa�s������� 3�N�߿���(�:� ̿]�oρϔ�'�9�ʯ �������$���H�Y� k�}ߐ���+�ƿ���� ��� ϻ�D�U�g�y� �Ϟ�1���������� ߭�@���c�u����� ��5�P������� <���_q���)�;� �������J� [m����(:L���/u�<s10712 ��^/�p/�/t7����'/2�/�/�/�/.�/0( �/]?o?�?&�4$ P?�?�?O�r�?+-��?bOtO�Optp�disc 0=O2� 9OKO�O�O _v�tpconn 0 �O�O�O[_m__�/ �/-?�/�_�_�_?"? �_F?Woio{o�?�?3O �?�o�o�oOO�oB_ 	ew
�_�_7oR ���o�>o�a� s����o+8��oߏ� �����L]�o��� ��/��۟�����$���H�Y�k�}�����$SNPX_AS�G 2������� � R"%���Я  �?���PARAM� ���� W�	��PӤ��9Ө$�������OFT_KB_CFG  ӣ�����OPIN_SIMW  ���}����������RVNO�RDY_DO  �)�U���QST_P_DSBi��|ϐ�SR �� � &#�D�O��O�:�TOP_ON_ERRʿ��o��PTN ��ޢ��A��RI?NG_PRMy�ܲ�VCNT_GP �2��!���x 	���ϗ���#��G����VD��RP 1	��"�8Ѩ�*߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�}�z��������� ������
C@R dv������ 	*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?[?X?j?|?�?�?�? �?�?�?�?!OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLosopo�o �o�o�o�o�o�o  96HZl~�� ������ �2��D�V�`�PRG_CoOUNTJ���N{�ENB��}�M���L���_UPD 1}'�T  
k� �����"�K�F�X�j� ��������۟֟��� #��0�B�k�f�x��� ������ү������ C�>�P�b��������� ӿο����(�:� c�^�pςϫϦϸ��� ���� ��;�6�H�Z� ��~ߐߢ��������� �� �2�[�V�h�z� ������������
� 3�.�@�R�{�v����� ��������* SN`r���t��_INFO 1��Ҁ� 	� ��3?�ڪK@T�?~ſc�8:�$�/�A8����e���8��8m��f��� DC@8�D��DH  �3��´���YSDEBUG���퀍dՉ�SP_�PASS��B?~+LOG �]��  � ���  �с�UD1:\;$�<"_MPCA-셽/�/��x!�/ 쁝&SAV D)����d!|"�%�(SV��+TEM_TIM�E 1D'�� 0Ҁ�΄u4�?�.�TMEMBK  	�сd d/�?�?��<X|Ҁ� @�?C�O:OJLHOmOzI�J��@p1�O�O�O�O"3 _�_$_6_H_Z_l_ � n_�_�_�_�_�_�_�_o"o\�e1oVohozo �o�o�o�o�o�o�o
 .@Rdv���O5SK�0�8���?����F:� j��O%O΄AJ� p0p��3�\O����(�O!��Oя�����Ov4� � �j�9�G�f�x���~_!����ӟ���	��� $�C�7o g�y���������ӯ� ��	��-�?�Q�c�u�����������T1SVGUNSPD%%� '%��2M�ODE_LIM #a9"ܴ2�	�� D-۵ASK_?OPTION �9�!F�_DI ENB  U�%f��BC2_GRP 2!�u#o2��XB���C����ԼBCCF�G #��*< ��`ߐI� 4�Y��jߣߎ��߲� ��������E�0�i� T��x��������� ���/��S�>�w�����t���u�����c� ��	B-f�.� �4[ ������ � 02Dzh �������/ 
/@/./d/R/�/v/�/ �/�/�/�(���/?&? 8?J?�/n?\?~?�?�? �?�?�?�?O�?4O"O XOFOhOjO|O�O�O�O �O�O�O__._T_B_ x_f_�_�_�_�_�_�_ �_oo>o�/Voho�o �o�o(o�o�o�o�o (:Lp^�� ������ �6� $�Z�H�~�l������� ؏Ə��� ��0�2� D�z�h���To��ȟ� ��
���.��>�d�R� ������z�Я����� ��(�*�<�r�`��� ������޿̿��� 8�&�\�Jπ�nϐϒ� �������ϴ��(�F� X�j��ώ�|ߞ��߲� �������0��T�B� x�f���������� ����>�,�N�t�b� ���������������� :(^�v�� ��H���$ HZl:�~�� �����2/ /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?P?R? d?�?�?�?t�?�?O O*O�?NO<O^O�OrO �O�O�O�O�O�O__ 8_&_H_J_\_�_�_�_ �_�_�_�_�_o4o"o XoFo|ojo�o�o�o�o �o�o�o�?6Hf x���������v&��$TBC�SG_GRP 2�$�u� � �&� 
 ?�  Q�c�M��� q��������ˏ���*�1�&8�d,� �F�?&�	 H�CA��>�f�fb�N��CS��B�I�����V��3�3��n�C
��ԝB]�����&h���Blt�\ԟ�A���L��;���.�C�{����������G�w�CHd��k�LƯ��C�����@�� I��-���
�X�u�@��R�����̻�����	�V3.00I�	Omt7���*�� �%��ֶ:�H?�� &�H�� qN� �O�  ������ ϏϘ�*�J�21�'8��Ϥ�C�FG )�u�B� E������d�#��#�I�W� �pW�}�hߡߌ��߰� �������
�C�.�g� R��v�������� 	���-��Q�<�u�`� r�����������I� cp"4��gRw ������	 -?�cN�r� �&������/ </*/`/N/�/r/�/�/ �/�/�/?�/&??J? 8?Z?\?n?�?�?�?�? �?�?O�? OFO4OjO XO�O�O`�O�OtO�O _�O0__T_B_x_f_ �_�_�_�_�_�_�_�_ ,ooPoboto�o@o�o �o�o�o�o�o�o( L:p^���� ���� �6�$�F� H�Z���~�����؏Ə ����2��OJ�\�n� ������������ �
�@�R�d�v�4��� ������ί����ү (�N�<�r�`������� ��ʿ̿޿��8�&� \�Jπ�nϐ϶Ϥ��� ������"��2�4�F� |�jߠߎ����߀���  �߼�B�0�f�T�� x����������� �>�,�b�P������� ��v�������: (^L�p��� �� �$H6 lZ|����� �/�/ /2/h/�� �/�/�/N/�/�/�/
? �/.??R?@?v?�?�? �?j?�?�?�?�?O*O <ONOOO�OrO�O�O �O�O�O�O _&__J_ 8_n_\_�_�_�_�_�_ �_�_o�_4o"oXoFo ho�o|o�o�o�o�o�o �/$6�/�oxf �������� ,�>���t�b����� ��Ώ��򏬏��&� (�:�p�^��������� ܟʟ�� �6�$�Z� H�~�l�������دƯ ��� ��D�2�T�z� h���Jȿڿ���� ��
�@�.�d�Rψ�v� �Ͼ����Ϡ����� �*�`�r߄ߖ�Pߺ� �����������&� \�J��n������ ������"��F�4�j� X�z�|����������� ��0B�Zl~ (������� ,Pbt�D�������   # &0/"��$TBJOP_�GRP 2*���  K?�&	H"O#,V,����x�� =k% � �< ��� �$ @� g"	 �CA����&��SC��q_%g!�"!G��"�Q��/� .{�2^�R=��CS�?���?�&0L��B�  B<�'??J7�/��/?(��6}? �?(�à5;���v 6�*?<?�;B�~�7C�  D�!�,0��B�0OK�:�Z�Bl  �@pB@�ff?�/�
CH�0��?gOO  A�zG�2jG��&�5333�O�K;g��|A�!@J@_�ffC�Z0zjO�Oz@���U�O�$�#�
0R�E1_CV;�xCsQ@���@&ff@���O�_tF�X_�$:�H�RJ=q�_�8AP�:�t-�Q?�33@�@@�Oo�_ ,i$oZGLo6oDoro�o ~o8o�o�o�o�o3 �oRlVd���V4�&b x�%	�V3.00m#'mt7A@�s*�l$�!�'� E���qE���E��]\E�HF�P=F�{F*�HfF@D�FW��3Fp?F��MF���F��MF��F��şF��F��=F���G��G.8�C�W�RD3l)D���E"��E�x�
E��E��,)FdRF�BFHFn� F���F��MF��ɽF�,
G�lGg!G�)�G=��G�S5�GiĈ;^M@;�o�|# 2 dXz&/��5&"�?��PYO�WOE#ESTPAR�S  (a E#H�Rw�ABLE 1�-V) @�#DR�7� � �R�R��R�'#!R�	R�
�R�R���!R��R�R���RDI��`!��ԟ���
�r�Oz���������H̯ޮ��Sx�^# <� ����ÿտ����� /�A�S�e�wωϛϭ� ��������;-w�{�_" ��6��1�C�U����%�7�I�[����NUoM  �`!� $  ��m���_CFG .�����BH IMEBF_TT}���^#��G�GVERk�H�]�G��R 1/�� 8I�" �� �A�  ��������� ��� �2�D�V�h�z� ������������/
 e@Rhv�� �����* <N`r���� ��'///]/8/J/ `/n/�/�/�/�/r���_��t�@~�t�M�I_CHANS� �~� !3DBGLV�LS�~�s�$0ET�HERAD ?*��w0�"��/�/�?�?l�$0ROUT6q�!�!�4�?~�<SNMASKl8|~�}1255.2E��s0OBOTO�st�OOLOFS_DI}���%V9ORQCTRL 0���#��MT�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo&l�OIo8o�moq�PE_DET�AIJ8�JPGL_�CONFIG �6�ᄀ/c�ell/$CID?$/grp1qo�o �o/壀�?Z l~���C�� �� �2��V�h�z� ������?�Q����
� �.�@�Ϗd�v����� ����M������*� <�˟ݟr���������̯@�}a���&�8�@J�\���^o��c��`� ��˿ݿ���Z�7� I�[�m�ϑ� ϵ��� �������!߰�E�W� i�{ߍߟ�.������� �����A�S�e�w� ����<�������� �+���O�a�s����� ��8�������' 9��]o���� F���#5� Yk}�����`��User �View �i}}�1234567890�//,/>/P/�X$� �cx/���2 �U�/�/�/�/??s/�/�3�/b?t?�?@�?�?�??�?�.4Q? O(O:OLO^OpO�?�O�.5O�O�O�O __$_�OE_�.6�O~_�_��_�_�_�_7_�_�.7 m_2oDoVohozo�o�_�o�.8!o�o�o
�.@�oagr �lCamera��o����� �ޢE�*�<�N���h�z��������I  �v�)��$�6�H� Z�l����������؟@���� �2�Y��v P9ɟ~�������Ưد ���� �k�D�V�h� z�����E�W�I5�� ��� �2�D��h�z� ��׿����������
� ��W�ދ��X�j�|ߎ� �߲�Y�������E�� 0�B�T�f�x�߁ulY ���������
���� @�R�d���������� ������W� iy�.@ Rdv�/���� �*<N�� W��i������ ��/*/</�`/r/@�/�/�/�/as9F/ �/??1?C?U?�f? �?�?D/�?�?�?�?	O(O-O�j	�u0�?hO zO�O�O�O�Oi?�O�O 
_�?._@_R_d_v_�_ /OAO�p�{,_�_�_o o)o;o�O_oqo�o�_ �o�o�o�o�o�_�u ���oM_q��� No���:�%�7� I�[�m�NEa���� ˏݏ����7�I� [����������ǟٟ ����ͻp�%�7�I�[� m��&�����ǯ�� ���!�3�E�쟒�9� ܯ������ǿٿ뿒� �!�3�~�W�i�{ύ� �ϱ�X�����H���� !�3�E�W���{ߍߟ� ��������������  ��L�^�p� ����������� ��   "�*�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������//�*/</N/`/r/�/� � 
��(  �>@�( 	 �/�/ �/�/�/? ?6?$?F? H?Z?�?~?�?�?�?�*2� �l�O/O AO��eOwO�O�O�O�O ��O�O�O_TO1_C_ U_g_y_�_�O�_�_�_ _�_	oo-o?oQo�_ uo�o�o�_�o�o�o�o ^opoM_q�o ������6� %�7�~[�m������ ���ُ���D�!�3� E�W�i�{�ԏ��ß ՟�����/�A�S� ��w�����⟿�ѯ� ����`�=�O�a��� ��������Ϳ߿&�8� �'�9π�]�oρϓ� �Ϸ���������F�#� 5�G�Y�k�}��ϡ߳� ���������1�C� �ߜ�y��������� ����	��b�?�Q�c� �������������(� )p�M_q�p�����0@ �������� ���#frh:\t�pgl\robo�ts\m10ia�4_7l.xml �Xj|����0���.��/1/ C/U/g/y/�/�/�/�/ �/�/�//?-???Q? c?u?�?�?�?�?�?�? �?
?O)O;OMO_OqO �O�O�O�O�O�O�OO  _%_7_I_[_m__�_ �_�_�_�_�__�_!o 3oEoWoio{o�o�o�o �o�o�o�_�o/A Sew����� ��o��+�=�O�a� s���������͏ߏ�:I ��<<  ?��4��,�N�|�b� ������ʟ�Ο��� 0��8�f�L�~�����Д��������(��$TPGL_OUTPUT 9������  $�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ������$����2345678901�� � �2�D�V�^����� �ߗߩ߻�����w���@�'�9�K�]���}g� ��������o��� �1�C�U�g���u��� ��������}���- ?Qc����� ����);M _q	���� ���%/7/I/[/m/ //�/�/�/�/�/�/ �/?3?E?W?i?{?? %?�?�?�?�?�?O�? OAOSOeOwO�O!O�O��O�O�O�O_�O� $$Ӣ��OW =_o_a_�_�_�_�_�_ �_�_�_#ooGo9oko ]o�o�o�o�o�o�o�o@�oC5g}���������}@���"�� ( 	 iW�E�{�i� ����Ï��ӏՏ�� �A�/�e�S���w��� �����џ���+���;�=�O���s����Ƹ  <<\ ޯ�)�ͯ�)��M� _���ʯ����<���ؿ ��Ŀ� �~�$�V�� BόϞ�x�����2ϼ� 
ߤ���@�R�,�v߈� ��p߾���j������ �<�߬�r���� �������`�&�8� ��$�n�H�Z������ ��������"4X j��R��L�� ��|Tf  ��v��0B/ /�&/P/*/</�/�/ ��/�/h/�/??�/ :?L?�/4?�??n?�? �?�?�? O^?�?6OHO �?lO~OXO�O�OO$O �O�O�O_2___h_ z_�O�_�_J_�_�_�_��_o.o��)WG?L1.XML�cm��$TPOFF_�LIM Š�p����qfN_S]Vy`  �t�j�P_MON :����d�p�p2�miSTRTCHK' ;���f~tb�VTCOMPAT��h*q�fVWVAR� <�mMx�d K e�p�b�ua_DEFPR�OG %�i%�|�rd_DISP�LAY�`�n�rIN�ST_MSK  ��| �zINU�SER �tLCK�)��{QUICKM�ENM��tSCRE�l���+rtpsc�t)������b���_��STz�iR�ACE_CFG �=�iMt�`	�nt
?��HNL� 2>�z���T{  zr@�R�d�v����������К�ITEM �2?,� �%$�12345678�90�%�  =<��C�U�]�  !c�k�wp'���ns� ѯ5����k������ j�ů��鯕���A�1� C�U�o�y�󿝿I�o� ��忥�	��-ϧ�Q� ��#�5ߙ�A߽����� e߳������M���q� ��L��g��ߋ��� ��%�w� �[���+� Q�c���o�������� 3���{�;���� ��G_����/� Se.�I�m ���=�a /3/������ k//�/�/�/]/?�/ �/�/?�/u?�?�?? �?5?G?Y?�?+O�?OO aO�?mO�?�?�OO�O CO__yO+_�O�Ox_ �O�_�O�_�_�_?_�_ c_u_�_o�_Wo}o�o �_�oo)o;o�o�oqo 1C�oO�o�o� �%��[���Z��S�@��_�ψ  ے_� 8����y
 Ï��Џ���UD1:�\���q�R_G�RP 1A �?� 	 @�pe� w�a���������ߟ͞����ّ�>�)�<b�M�?�  }��� y�����ӯ������ 	��Q�?�u�c�����0����Ϳ�	-����o�SCB 2B{� h�e�wωπ�ϭϿ�������e�U�TORIAL �C{��@�j�V_C�ONFIG D�{���������O�OUTPUT E{���������� �%�7�I�[�m��� ������������ %�7�I�[�m������ ����������!3 EWi{���� ����/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/��/? ?'?9?K?]?o?�?�? �?�?�?�/�?�?O#O 5OGOYOkO}O�O�O�O �O�O�?�O__1_C_ U_g_y_�_�_�_�_�_ �O�_	oo-o?oQoco uo�o�o�o�o�o�_�o );M_q� �����yߋ��� �-�?�Q�c�u����� ����Ϗ���o�)� ;�M�_�q��������� ˟ݟ� ��%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� 
��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ���1CUgy �������	 -?Qcu��������/�x���$/6/ !/ a/��/�/�/�/�/�/ �/??'?9?K?]? �?�?�?�?�?�?�?�? O#O5OGOYOkO|?�O �O�O�O�O�O�O__ 1_C_U_g_xO�_�_�_ �_�_�_�_	oo-o?o Qocot_�o�o�o�o�o �o�o);M_ q�o������ ��%�7�I�[�m�~ ������Ǐُ���� !�3�E�W�i�z����� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o��~��$TX_SCREEN 1F8%�  �}�~���������
�����m&}/FR�/testeIH�M.stm K � g����g ��T�(��'����Kgӈ�o�ɯ}m%S�(,���t�m)����aӛ�}�tг��v=,ѿTELA1j��?��'܈�^֯� ��
��.�@�R�-�?� h����������f� x�%�7�I�[�m���� �����������! ����<i{��� �:L�/A S�w����� ��l~/=/O/a/�s/�/�//��UAL�RM_MSG ?5����� �/�� �/�/)??M?@?q?d? v?�?�?�?�?�?�?O~�%SEV  �-�EF�"ECFG� H���� � ��@�  A�uA   Bȁ�
 O���ŨO�O�O �O�O__&_8_J_\_�jWQAGRP 2I�[K 0��	 ��O�_� I_BBL�_NOTE J�[JT���l������g@�RD_EFPRO� %�+ (%O.o��o Uo@oyodo�o�o�o�o��o�o�o?�\F�KEYDATA �1K�ɞPp jG�� h_��`�P����u,(J ����J�1�n�U��� ����ȏ������"� 	�F�X�?�|�c����� ��֟������0��T��~��d������� ��ӯ寈�y�� �2� D�V�h���������¿ Կ�u�
��.�@�R� d�v�ϚϬϾ����� �σ��*�<�N�`�r� ߖߨߺ�������� ��&�8�J�\�n��� ������������"� 4�F�X�j�|������ ����������0B Tfx���� ���>Pb t��o����� //:/L/^/p/�/ �/�/5/�/�/�/ ?? $?�/H?Z?l?~?�?�? 1?�?�?�?�?O O2O �?VOhOzO�O�O�O?O �O�O�O
__._�OR_ d_v_�_�_�_�_M_�_ �_oo*o<o�_`oro �o�o�o�oIo�o�o &8J�on�� ���W���"� 4�F��j�|�������hď֏�܋�������)��K�]�7�,I���A� ����֟�ϟ��0� B�)�f�M��������� �����ݯ��>�%� b�t�[������ο� ���(�:�L�[�p� �ϔϦϸ�����k� � �$�6�H�Z���~ߐ� �ߴ�����g���� � 2�D�V�h��ߌ��� ������u�
��.�@� R�d������������ ������*<N` r������ &8J\n� ������� "/4/F/X/j/|//�/ �/�/�/�/�/?�0? B?T?f?x?�?�/�?�? �?�?�?OO�?>OPO bOtO�O�O'O�O�O�O �O__�O:_L_^_p_ �_�_�_5_�_�_�_ o o$o�_HoZolo~o�o �o1o�o�o�o�o  2�oVhz��� ?���
��.�� R�d�v���������M� ����*�<�ˏ`� r���������I�ޟ�@��&�8�J�!0L���!0����u�����q���ͯ��, ������"�	�F�X�?� |�c�������ֿ���� ��0��T�f�Mϊ� qϮϕ���������� ,�>�?b�t߆ߘߪ� ��˟������(�:� L���p������� Y��� ��$�6�H��� l�~�����������g� �� 2DV��z �����c�
 .@Rd��� ����q//*/ </N/`/��/�/�/�/ �/�/�//?&?8?J? \?n?�/�?�?�?�?�? �?{?O"O4OFOXOjO |OSߠO�O�O�O�O�O O_0_B_T_f_x_�_ _�_�_�_�_�_o�_ ,o>oPoboto�oo�o �o�o�o�o�o: L^p��#�� �� ���6�H�Z� l�~�����1�Ə؏� ��� ���D�V�h�z� ����-�ԟ���
� �.���R�d�v����� ��;�Я�����*� ��N�`�r���������ڑ@����@������	��+�=��,)�n�!ߒ�y� ���ϯ������"�	� F�-�j�|�cߠ߇��� �߽�������B�T� ;�x�_���O���� ����,�;�P�b�t� ��������K����� (:��^p�� ��G�� $ 6H�l~��� �U��/ /2/D/ �h/z/�/�/�/�/�/ c/�/
??.?@?R?�/ v?�?�?�?�?�?_?�? OO*O<ONO`O�?�O �O�O�O�O�OmO__ &_8_J_\_�O�_�_�_ �_�_�_�_��o"o4o FoXojoq_�o�o�o�o �o�o�o�o0BT fx����� ���,�>�P�b�t� �������Ώ���� ��(�:�L�^�p���� ����ʟܟ� ���� 6�H�Z�l�~������ Ưد������2�D� V�h�z�����-�¿Կ ���
�ϫ�@�R�d� vψϚ�)Ͼ����������*�`,��>`���U�g� y�Qߛ߭߇�,���� �����&�8��\�C� ���y��������� ���4�F�-�j�Q��� u����������� �_BTfx���� ����,� Pbt���9� ��//(/�L/^/ p/�/�/�/�/G/�/�/  ??$?6?�/Z?l?~? �?�?�?C?�?�?�?O  O2ODO�?hOzO�O�O �O�OQO�O�O
__._ @_�Od_v_�_�_�_�_ �___�_oo*o<oNo �_ro�o�o�o�o�o[o �o&8J\3 �������o� �"�4�F�X�j���� ����ď֏�w��� 0�B�T�f��������� ��ҟ������,�>� P�b�t��������ί �򯁯�(�:�L�^� p��������ʿܿ�  Ϗ�$�6�H�Z�l�~� Ϣϴ���������� ��2�D�V�h�zߌ�� ����������
��.�@�R�d�v���qp����qp���������������,	N�r�Y����� ����������& J\C�g��� ����"4X ?|�m���� �/�0/B/T/f/x/ �/�/+/�/�/�/�/? ?�/>?P?b?t?�?�? '?�?�?�?�?OO(O �?LO^OpO�O�O�O5O �O�O�O __$_�OH_ Z_l_~_�_�_�_C_�_ �_�_o o2o�_Voho zo�o�o�o?o�o�o�o 
.@�odv� ���M���� *�<��`�r������� ��̏�����&�8� J�Q�n���������ȟ ڟi����"�4�F�X� �|�������į֯e� ����0�B�T�f��� ��������ҿ�s�� �,�>�P�b��Ϙ� �ϼ������ρ��(� :�L�^�p��ϔߦ߸� ������}��$�6�H� Z�l�~�������� ����� �2�D�V�h� z�	��������������
������5GY1{�g,y�q� ��<#`r Y�}����� /&//J/1/n/U/�/ �/�/�/�/�/�/ݏ"? 4?F?X?j?|?���?�? �?�?�?�?O�?0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�_�_'_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  $�oHZl~�� 1����� �� D�V�h�z�������?� ԏ���
��.���R� d�v�������;�П� ����*�<�?`�r� ����������ޯ�� �&�8�J�ٯn����� ����ȿW�����"� 4�F�տj�|ώϠϲ� ����e�����0�B� T���xߊߜ߮����� a�����,�>�P�b� �߆��������o� ��(�:�L�^���� ������������}� $6HZl���� ����y 2�DVhzQ�|}�Q�����@������,�/ ./�/R/9/v/�/o/�/ �/�/�/�/?�/*?<? #?`?G?�?�?}?�?�? �?�?OO�?8OO\O nOM��O�O�O�O�O�O �_"_4_F_X_j_|_ _�_�_�_�_�_�_�_ o0oBoTofoxoo�o �o�o�o�o�o�o, >Pbt��� �����(�:�L� ^�p�����#���ʏ܏ � ����6�H�Z�l� ~������Ɵ؟��� � ���D�V�h�z��� ��-�¯ԯ���
�� ��@�R�d�v������� �Oп�����*�1� N�`�rτϖϨϺ�I� ������&�8���\� n߀ߒߤ߶�E����� ���"�4�F���j�|� ������S������ �0�B���f�x����� ������a���, >P��t���� �]�(:L ^������� k //$/6/H/Z/� ~/�/�/�/�/�/�/����+������?'?9=?[?m?G6,YO�?QO�?�?�? �?�?OO@ORO9OvO ]O�O�O�O�O�O�O_ �O*__N_5_r_�_k_ �_�_�_�_��oo&o 8oJo\ok/�o�o�o�o �o�o�o{o"4F Xj�o����� �w��0�B�T�f� x��������ҏ��� ���,�>�P�b�t�� ������Ο������ (�:�L�^�p������ ��ʯܯ� ���$�6� H�Z�l�~������ƿ ؿ���ϝ�2�D�V� h�zό�ϰ������� ��
���_@�R�d�v� �ߚߡϾ�������� �*��N�`�r��� ��7���������&� ��J�\�n��������� E�������"4�� Xj|���A� ��0B�f x����O�� //,/>/�b/t/�/ �/�/�/�/]/�/?? (?:?L?�/p?�?�?�? �?�?Y?�? OO$O6O�HOZO�$UI_I�NUSER  ����{A?�  [O_O�_MENHIST� 1L{E  ( �@���'/SOFT�PART/GEN�LINK?cur�rent=men�upage,71�,1�O__0_B_ �O�O,74�O�_�_ �_�_S_e_�A3|_o�#o5oGo�2)�_�_8 �@o�o�o�o�o�_po,37o,>Pr�1(�oj^955	������ov�q8 �"�4�F�X�c��r�36�����ˏݏ  ���0�A���� "�4�F�X�j� ���� ����şן�x��� 1�C�U�g��������� ��ӯ������-�?� Q�c�u��������Ͽ �󿂿�)�;�M�_� qσ�ϧϹ������� ��%�7�I�[�m�� �ߔϵ���������� ��3�E�W�i�{��� �������������� A�S�e�w�����*��� ��������=O as���8�� �'�0]o �������� /#/5/�Y/k/}/�/ �/�/B/�/�/�/?? 1?C?�/g?y?�?�?�? �?P?�?�?	OO-O?O �?POuO�O�O�O�O�O ^O�O__)_;_M_8 �O�_�_�_�_�_�_�O oo%o7oIo[o�_o �o�o�o�o�o�ozo !3EWi�o�� ����v��/� A�S�e�w�������� я������+�=�O��a�s�^[�$UI_�PANEDATA 1N������  	��}/FR/t�esteIHM.�stm Ñ?_w�idth=0&_�height=1�0Ԑdevice�=TP&_lin�es=3Ԑcol�umns=4Ԑf�onܐ4&_page=doub��1��\V)pri9m#�L�  }O�s�`��������ͯ )ϯ �گ���;�M�4�q� X�������˿������%�\V�� �E�  w���]�d/frh/�cgtp/flex�ȟڟ2����y2/�-�dual�� ��_��"�4�F�X�j� ώ�u߲��߫����� ���B�)�f�M�ﰜ����3� G��������*�<�N� `�����Ϩ������� ��i�&8\C ��y�������4Xj=�  ����������� � /S$/��H/Z/l/ ~/�/�/	/�/�/�/�/ �/ ?2??V?=?z?a? �?�?�?�?�?�?
O} �@OROdOvO�O�O�? �O1/�O�O__*_<_ N_�Or_Y_�_}_�_�_ �_�_�_o&ooJo1o no�ogo�oO)O�o�o �o"4�oXj�O ������O� �0�B�)�f�M����� ���������ݏ�� >��o�o��������� Ο��3��w(�:�L� ^�p���韦�����ܯ ï ����6��Z�A� ~���w�����ؿ�]� o� �2�D�V�h�z�Ϳ �����������
�� .ߕ�R�9�v�]ߚ߬� ���߷������*��@N�`�G����	����@���������"�)�� G���6�s��������� ��4�������K 2oV���������#������$UI_POST�YPE  ��� 	 �/�UQUICK�MEN  d�s�WRESTO�RE 1O��  ���� /#���m +/T/f/x/�/�/?/�/ �/�/�/?�/,?>?P? b?t?/�?�?�??�? �?OO(O�?LO^OpO �O�O�OIO�O�O�O _ _�?_1_C_�O~_�_ �_�_�_i_�_�_o o 2o�_Vohozo�o�oI_ So�o�oAo�o.@ Rd����� s���*�<��oI� [�m������̏ޏ�� ���&�8�J�\�n���������ȟڟ�SC�RE�?��u1sc�uU2�3�4�5��6�7�8��T;AT`� ��MUSER�����Sks���3��4��U5��6��7��8���UNDO_CFG� Pd����UP�DX�����None���_I�NFO 1Q�<��0%��W��� E���i��������� տ���:�L�/�pς��eϦύ)�OFFS�ET Td@� ��{������	��-� Z�Q�cߐ߇ߙ��ϝ� ������ ��)�V�M�_�q�۹�����
����t��)�WOR/K U4������A�S��ψ�UFRAME  ���&��RTOL_ABRqT��$���ENB��~��GRP 1V���Cz  A� ��+=Oa s�����U����~��MSK  ��<���N��%4���%��)��_EVN������>�2W���
 h��U�EV��!td:�\event_u�ser\-�C7ȍ��}�F��SP���spotw�eld�!C6 ����!� Z/�/:'�H/~/l/�/ �/�/�/-?�/Q?�/?  ?�?D?�?h?z?�?O �?)O�?�?OqO`O�O @ORO�OvO�O_�O�O@7_�O[__Z]W+�32X����8V_�_�_ �_�_o�_,o>o obotoOo�o�o�o�o �o�o�o:L'�p�]����$�VARS_CON�FI�Y�� FP�{���|CCRG��\��>�{��t�D� BH� p,k�a�C�� ��}��?���C,&Q=��mͩ�A �MR;2b���	}��	��@�%1: �SC130EF2� *����{�����,X� �5}������A@k�C�F� 	w�Q�[���|��� �������T�����\�ϟ �\� B���;�e�@�ǟ `�����S�����̯�� �ۯ�&�}��\�G��Y���E���ȿ�TCC�c
�������M�pGF�pgd���-�2345?6789017�?��ׁ$���4�v�N m�� ��϶�BW������i�}�:�o=LA�څ�6�@�6�Ϳ�Z���i�7����(�� W���-�]�X�jĈߚ� �ϳϹ��������� %�7�I�r�m�ߨ�� �����������8�3� E�W������}����� ��������/�A�S�xe�w��MODE���t �RSLTg e�|k�%"z� ���;�1��d���`��SELEC���c��	IA_[WO�Pf ��� W,		�������G�P ������RTSYONCSE� ��$��	#WINURL 3?*ـ�;\/�n/�/�/�/�/�uISIONTMOU����A# ��%�g�Sۣ�SۥP��� FR:\~�#\DATA\�/� �� MC�6LOG?   oUD16EX@?�\�' B@ ���2T1���?T1�?�?����� n6  ���GV<�2\� -��5��   ��Z�@�U058TRAIN�j?��*B{Rd_Cp���F#`{2��'$�"��h#� ( �kI�Mw��O�O�O�O �O1__U_C_]_g_y_p�_�_�_�(STA� 	i��@�?o0oI:q$obo�%_GE��j#��~@ �
�\��btgHOMI}N�kSۮ��`��2,,��CWǖ�BveJMPERR� 2l#�
   QoI:��"�4Fw j|����������&%S_g0R�E�m�^۴LEXzdn�1-eho�VMPHASE � �e׃BޱO�FF _ENB { �$VP2�$_oSۯ��x�c
 C;�@ �@�;���?s33'D*AA��]� ��0ޱ
�`r}�XC��܅�ๆ\A-۟E  ������#�5����� ��������}������ ����c�X���A��� ��ϯ�+��߿�� M�B�q���xϊϹ��� Ϸ�������7�I�;� m�b�)ߣ�Eߓߡ߳� ����3���W�L�{� ���ߑ��������� �/�$�6�e�W���c� y������������ ��O���?M_q�� �����'9� =7Is���� ��/m/%/3/�E/s�TD_FIL�TE�`s�k �x2�`����/�/�/ �/�/	??-???Q?�6 �/~?�?�?�?�?�?�?��?O OoiSHIF�TMENU 1t}<5�%5�~O)� \O�O�O�O�O�O�O�O '_�O_6_o_F_X_�_�|_�_�_�_	LIVE/SNAP�Svsfliv����_�z`ION� ҀU
`bmenu&o+o�_�o�oV"<Ej�uz��4IMO��v���zq�WAI�TDINEND � �ec��b�fOK�وOUT�hS�DyTIMdu��o|G�}#�{C��zb�z�xREL1E��ڋxTM�{�d{��c_ACT`�و��x_DATA' wz���%�oď<5Fx�RDIS
`E���$XVR�a�x�n�$ZABC_GRP 1yz���� ,�2�̏.MZD��CSC%H�`z���aP@�h�@�IP�b{�'���şן�[�M�PCF_G 1|
'���0�r�8���� �}'��p�s�� 	(���  <�l0  �����3_=?� ? 4M���������3�DC�@8D��DH��1w��Dq >�Nnl��`��?Nng5��z��� ��ïկ�����o�p��w���� /�?�3��´ſ׾ ĸ��	��1�?�i���'��0?�Q���	��`~����_CY�LIND~!�� Р ,(  *.�?ݧ+�h�O���s� �������� (�	�x�-��&�c�� ��������j�P�� ��)��~�_�q��� �s2�'��� �&� ���������&���I��cA���S�PHERE 2��������� �A�T/A��e ������/ N`=/�a/H/Z/�/`��/�/�/�ZZ� ��f