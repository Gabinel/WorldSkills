��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@  &��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	4SU�SRVI 1  < `�R*�R�n�QPRI�m� �t1�PTRIP�"m��$$CLASP ����a��R2��R `\ SI�	g�  0�aIRTs1	o`�'2 L1�L1���R	 ,��?���a1`��b�d~a��a��� �  y����
 ��a��o�o1CU  �oz�����c �
��.�@�R��v� ��������Џ�q�� �*�<�N�`���� ����̟ޟm���&� 8�J�\�n��������� ȯگ�{��"�4�F� X�j���������Ŀֿ����`TPTX�����/�`� sȄ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ��� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F�X���|��������������a�f�oC ($ p�-����T�?�x���a�a��c���c����l��c�g�e�a�a�dh��a2�h�\�Ph�����������`���`  ����f ep���h#h�F�bc �Xc�B 1)hR� \ _��� REG V�ED]���wh�olemod.h�tm�	singl�	doub �trip8browsQ�� ���u���/�/@/���dev.sl�/3� 1�,	t�/_�/;/ i/??/?�/S?e?w?8�?�?�?� ��? �?OO%O7OIO[OmO O�E2P�?�O�O�O�O �O_�E�	�?�?;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo oM'�o�o�o�o�o�o +=Oas� ��������? >�P�b�t��������� Ώ���O�����L� ^�_'_�������ş �����6�1�C�U� ~�y�����Ư��ӯ�o ���-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�-��Ϭ� ����������*�<� 7�`�r�A�Sߨߺ�q� ��i�����!�J�E� W�i��������� ����"��/���O�I� w��������������� +=Oas� ������, >Pbt���߼ ���//����� ^/Y/k/}/�/�/�/�/ �/�/�/?6?1?C?U? ~?y?�?Y��?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _�R_d_v_�_�_�_ �_�_�_�_�o*o�_�o`oro�j�$UI�_TOPMENU� 1K`�aR 
d�a�*Q)*defa�ult5_]*�level0 * [	 �o�0��o'rtpio�[23]�8tpst[1[x)w9��o	�=h58E�01_l.png���6menu5�y�p�13�z��zb	�4���q��]� ��������̏ޏ)Rr����+�=�O�a����prim=�pa�ge,1422,1h�����şן����1�C�U�g����|�class,5�p�����ɯۯ�����13��*�<�N�`�4r���|�53�������ҿ�����|�8 ��1�C�U�g�y�����@����������"Y�` �a�o/��m!ηq�Y���avtyl}Tfqm�f[0nl�	��c�[164[w��59`[x�qG�y��tC8�|�29��o�%�1�� �{��m��!����� 0�B���f�x���������o���80�� '9K~���2P� ����\�� '9K����� �������1��/�$/6/H/Z/U�|�ainedi'ߑ/�/�/�/�/P�con�fig=sing�le&|�wintp���/$?6?H?Z?	��ߐ??ٷ�gl[57�ٳq��?�;gp�0	8�ݲ07I�?F��F2JO[6�:�?)O��O�x �� �4s�x�O���$��`� o�H_Z_l_~_�_�_Q� �_�_�_�_o o�_Do�Vohozo�o�o�o�!;^�$doub5o���13��&dual6�i38��,4�o&�o9�o�n�o�a8 ���Ao����(&�8��%3L=}!��o�b8@����������z���(�:��+:<T��i48,2o��b0{����ʟ {?�;�M�sc���;���s �� �}���e�u��X��@�F7L���`�OА�2�h�z�6e�u7 �����ｿϿ���̏�27��G�Y�k� }Ϗ��0�s������(���!�1�M� _�q߃ߕ�������� �����7�I�[�m� �������������!�����6(�]�o�`�������$��746�@����)�C�ߟ�T�	TPTX[G209�<Aw2IHJ���Bw1H�]H������02���A#��[Ttv `��O�L#_�0� \���5S[�treev'iew3v�3��~�?381,26M/ _/q/0�/�/�/�/�/ �/~/?%?7?I?[?m? �o/(��o5%���?�?&�?�A�?\1~��?8"2��eOwO�?�?( }�LEK��O�O_�O���8@�ONOa_s_�_��6 _d�E_�_�_�_oV� #_���_�Sooo�o�o B�o�o��oA�oq +=Oas� �o������� (�9���Q�x������� ��ҏ?����,�>� P�ߏt���������Ο ]�����(�:�L�^� ퟂ�������ʯܯk�  ��$�6�H�Z��l� ������ƿؿ�y��  �2�D�V�h����Ϟ� �������ϕo�o��o @ߧE�c�u߇ߙ߬� ������O����)�<� M�_�q���W����� ����&�8���\�n� ��������E������� "4��Xj|� ���S�� 0B�fx��� �O��//,/>/ P/�t/�/�/�/�/�/ ]/�/??(?:?L?�� ߂?1ߦ?���?�? �?�?O$O5OGO�?SO }O�O�O�O�O�O�O�O ��2_D_V_h_z_�_�_ �/�_�_�_�_
oo�_ @oRodovo�o�o)o�o �o�o�o*�oN `r���7�� ���&��J�\�n� ��������E�ڏ��� �"�4�ÏX�j�|��� ����a?s?蟗?�sO _/�A�S�e�w����� ����������,� =�O�a�#_������ο ��=��(�:�L�^� pς�Ϧϸ�������  ߏ�$�6�H�Z�l�~� ߐߴ���������� ��2�D�V�h�z��� ����������
���� @�R�d�v�����)����������ƚԔ�*default�%��*level8�ٯw���?� tpst[�1]�	�y�t?pio[23����u���J\�menu7_l.�png_|13���5�{�y4�u6���//'/ 9/K/]/���/�/�/�/ �/�/j/�/?#?5?G?�Y?k?�"prim�=|page,74,1p?�?�?�?�?��?�"�6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_�B_T_f_x_{?�218 �?�_�_�_�_�__B6o9oKo]ooo�o`��$UI_USE�RVIEW 1�֑֑R 
���o��o�o[m�o'9K ] �����l ���#�5��oB�T� f������ŏ׏鏌� ��1�C�U�g�
��� ������ӟ~����� v�?�Q�c�u���*��� ��ϯ�󯖯�)�;� M�_�
��~������ ݿ���%�ȿI�[� m�ϑ�4ϵ������� �Ϩ�
��.ߠ�i�{� �ߟ߱�T�������� �/���S�e�w��� Fߨ����>���+� =�O���s��������� ^�����'���� FX��|���� ��#5GY� }����p�� �h1/C/U/g/y// �/�/�/�/�/�/�/? -???Q?c?/p?�?�? ?�?�?�?OO�?;O MO_OqO�O&O�O�O�O �O�O�?�O_ _�OD_ m__�_�_�_X_�_�_ �_o!o�_EoWoio{o �o0h