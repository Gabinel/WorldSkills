��   �;�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_CPC�_T 4 $�COMMENT �$ENAB�LE  $M�ODJGRP_N�UMKL\  $UFRM\~] _VTX M ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�? �ELAY_T�IMJSPEED�_CTRLKOV�R_LIM? p JD� L��0�UTOO(i��O��&}S. � 8J\TC�u
!����\� �jY0  � ��CHG_SIZ��$AP!�E.�DIS�]$!B�C_+{#s%O#J�
p 	]$Jd#� �&s"��"{#�)�$�'�_S}EEXPAN#�N�iGSTAT�/ DFP_�BASE 5$0K$4!� .6K_V7>H73hJ- � }�\7AXS\UP�LW�7���
0c5r �< w?�?�?���?�?�//	7E�LEM/ T 1�&B.2NO�G]@�%CNHA�DF#� _$DATA)he0  PJ�@� 2 
&PN5 �� 1U*.n   _VSiSZHbRj0jR(�VyT(��R%S{TROBOT��X�SARo�U�V$CUR_��Rj�SETU4"	 ��bAISP_MGN��INP_ASS e#�PB!� `CiH�7�7`e�.fXc1�C�ONFIG_CH�K`E_PO* }dS/HRST�gM^#/e�OTHERRBTF�j_G]�R�dTv ��ku�c)&T1r
�0R HLH�d� 0  �lt<Ne'AVRF!YhH^t�5�1� �r�W�_A$Rdv�TPH/ (@G%Q�Q�Q3wwBOX/ 8�@ F!�F!�G �r{�z�TUIRi@ c ,�F�pER%@�2 $�p [L�_SF�!��ZN/ 0 �IF(@�p��Z_��0�_�0wu0 � @�Q7yv	
��~� �$$CL` ? �������Q��Q��VERS�ION���  0��IR�TUAL���' �2 �Q  ��p���&@>�m��P������P�������Ғd��Cz  0���� A���l���������Ɵ ۯ���� �2�D�F� h�}�����ԯſ��� ��
��.�@�R�d�f� �Ϛ�����п���ώ� �*�<�N�	�rχߖ� ��b��Ͼ�����&� 8�^�\�n߃��߶� ��������"�4�F� X�m�|�������� �����0�B�h�V x������������ ,>Pbw� ������// (:L�`/��/� ���/�??$/6/ H/Z/l/�?�/�?�/�/ �?�/�?O#O2?D?V? h?jO�?�O�?�?�?�O �O__.O@OROdOvO �O�_�_�O�O�_�O	o o�_<_N_`_r_-o�_ �o�_�_�o�_�o) 8oJo\o�o�o�o�2 �o�o��o�%�4F Xj|������� �����!�3�B�T�f� ��z�������ҏ��� ��/�>�P�b�t��� ������Ο������ +�=�L�^�p������ ��ʯܯ���'�9� H�Z�l�~����ϴ��� ؿ����#�5�G�V� h�zόώ߰������� ����1�C�R�d�v� �ߚ߬߮�������	� �-�?���`�r��� Q����������� ;M\�n��������� �V����"7I Xj|����� ���/E/W/f x���/��/�� /?,/A?S?b/t/�/ �/�/�?�/�?�/?O (?=OOOaOp?�?�?:O �O�?�O�? OO'_6O K_]_lO~O�O�O�O�_ �O�_�O_#o2_GoYo koz_�_�_�_�o�_�o �_
o@o1 Ugvo �o�o�o�o�o�� -�<Q�c���� ��u�����Ώ 8�*�_�q�������ʏ�ȏڋ�$DCSS�_CSC 2����Q  P����:�܉d
�k�.���R���v� ׯ����Я1���U� �y�<���`���ӿ�� �����޿?��c�u� 8ϙ�\Ͻπ��Ϥ�� ����;���_�"߃�F� ��j߷��ߠ����%� ��I��m�0���f���������GRPw 2�� ����	ҟS�>�w�b��� ������������ =(aL�p�� ���� K 6oZ�~��� ���/5/ /Y/D/ }/h/�/�/�/�/�/�/ ?�/
?C?.?g?R?�? �?�?z?�?�?�?�?O -OOQO<OuO�O�OdO �O�O�O�O_�O_;_ &___q_�_N_�_�_�_ �_�_�_�_%ooIo���_GSTAT 2���%��<� �� �+?�  ���?���6���5����3㴛�z���`A��Cj?��D+?���8`�<�e=.:~?�į䁴�aM2�ef^�a�a��`4���Z@�,�C��?����e�%��rdK>��i
�^l7���C.�r��`�g���s����C�? y��������?_�!���`�`4������+R�_cS���X������ �vC���<{�&Lp�Pq`p��du�c9�����A�y�`�DD�c�g9��`������Ts9�5���-5�x4��d�a��o�o�o y�� <�N���0�z���f��� Љ�i �-i��+k y  �.��&�H�v�\�~� �������ȟڟ��*� ��Z�l���x���|��� د���.��B��J� 0�B�d���x���ȿ�� ��������F�H�� �Ϻ�tϾ��Ϫ������͵���?��6<�R� �5���t��j�����P4�޿�5�@�K�C�"�D)���m<rEߎ?���c���1�~��c�ּ�m��b��C����m�Mq�Y�R?��� �gʿ�ٿY�e�������`C�� y���Q>��� �?r�;�q�<r�DN����e�њ�r�p������Ǹ��ӿ�C�ް�ڌ��-�����:�e��� �p��pK�&���@�M�C�ڑDB��� y<p]�?��)<�MJ����<pK9��/5��}�I�0�O� F�(�:�L��������� �� ����V�h��P� ��dϪ��������� ��F,^|bt ��j��8��< N(r�z���� �����,//4/ b/H/Z/|/�/�/�/�/ �/�"?T?X?j?D? �?�?z?���P�b�t� �ߘߪ߼�������� �(�:�L�^�p��O�? �?�?�?t_�_|?�_�_ �_�_�_o��/.o ? FodoJo\o~o�o�o�o �o�o�o�o2` ?���_���� � �odJ�xB�d� ��x���ȏ��Џ��� ���F�,�N�|�b�(� ����������*�<� �4_F_�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O_~�`�r��� ��"��.�X�2�D� �Ϡ�:����Ϝ��� � �����H�.�P�~�d� �ߴߚ߬����ߢ�,� >�p�*�t��`��� �� ������ �.�� 6�d�J�l��������� ����������Z�� F��|���п ⿈�������Я��� ��*�<�N�`�r��� ����/� ��/ �/��/�/�/�/*?<? ��$f?8~?�?�?�? �?�?�?�?O O2OPO 6OHOjO�O>�O�O? �O_"_�OF_X_N?�O �_�Oz_�_�_�_�_ o �_o6oo.oPo~odo �o�o�o`_�o(_�o, >btNl/~/$ 6HZl~��� ����/ /2/D/ �����VH�Z�P f���j�|�Ɵ؟r_�o ��o�8��0�R��� f�������ί�ү� �4��od�v���b��� ��������8��L� �8�f�L�nϜςϤ� �ϸ������ �"�P� 6�����Ŀ~����ߴ� ���������� ���,�>�P�b�t� ��������Ώ��R�4� F�X���������, bt�\ߞp� �����$ R8j�n��� v� //D�H/Z/4/ ~/�/���/��/�/ ?�/
?8??@?n?T? f?�?�?�?�?�?�?�/ .O`/OdOvOPO�O�O �O����\�n���� �����������"�4� F�X�j�|��_�O�O�O �O�o�o�O�o�o�o�o �o�/�?:ORp Vh������ �$�
��>�l�O�� ���o�����Џ�,� "p�V���N�p����� ��ԟ��ܟ
���$� R�8�Z���n�4�ʯ����� ���6�H�V���$DCSS_JP�C 2@�Q ( D=`��������P��ۿ ��������Y�(� g�Lϡ�p��ϔ��ϸ� ���1� ��g�6�H� Z߯�~��ߢ������ ��?�� �u�D�V�h� ���������)��� M��.�p���d�v��� ��������7[ *N�r��� ��!�/i8 �\������ �//�/"/w/F/�/ j/�/�/�/�/?�/�/ =???0?�?T?�?x? �?�?�?�?O�?�?8O ]O,O>O�ObOtO�O�O �O�O�O#_�OG__k_ :_L_�_p_�_�_�_�_��_��h�Sq�u�L �_Uooyo��dDo�o ho�o�o�o�o�o1 �oUy@Rd� ������?�� c�*���N���r����� 󏺏̏ޏ��M��q� 8���\�����ݟ��� ȟ%�����Y��F� ��j�ǯ��믲��֯ 3���W��e�B���f� x�����������A� �e�,ω�Pϭ�t��� �Ϫϼ��+���O�� s�:ߗ�^߻߂��ߦ� ������K��$�6� H��l�������� ��5���Y� �}�D�V� h������������� C
g.�R�v �������Q u<�`����/�&dMODE�L 23kx\��
 <�c (_  �z( �/g/y/�/�/�/�/�/ �/�/D??-?z?Q?c? u?�?�?�?�?�?�?.O OO)O;OMO_O�_�O Y/�O�O_�O�O<__ %_7_�_[_m_�_�_�_ �_�_�_�_8oo!ono EoWo�o{o�o�o�o�o �o�O�O�O�o|�o ew������ 0���+�=�O�a��� ����䏻�͏ߏ�� �b�9�K���3Es� ���m�۟����#� p�G�Y���}������� ůׯ$����Z�1�C� U�g�y���ؿ����� �������h��Q�c� �χϙ��Ͻ������ ��d�;�Mߚ�q߃� �ߧ߹�������N� %�7���1�C�q�� Y�����&����\�3� E�W�i�{��������� ����/A� ew������ �����=O�s �������/ P/'/9/�/]/o/�/�/ �/�/?�/�/:??#? 5?�?/]?o?�?�? �?O�?�?HOO1OCO �OgOyO�O�O�O�O�O �O�OD__-_z_Q_c_ �_�_�_�_�?
o�?�_ �_Ro)o;o�o_oqo�o �o�o�o�o�o< %7I[m��� ������!��_ ��oI�[�ȏ������ Տ�����/�|�S� e�����������џ� 0���f�=�O�a�s� ����m�������ѯ>� �'�t�K�]�o����� ���ɿۿ(����#� p�G�YϦ�}Ϗ��ϳ� ����$�������� 5�Gߴ�/ߝ߯����� ��2�	��h�?�Q�c� u����������� ��)�;�M���q��� ��k�}߫���*�� %7I[��� �����\3 E�i{���� /��F/����!/3/ �//�/�/�/�/�/? �/?T?+?=?O?�?s? �?�?�?�?O�?�?O PO'O9O�O]OoO�OW/ i/{/�O�O�O�O_^_ 5_G_�_k_}_�_�_�_ �_o�_�_Hoo1oCo Uogoyo�o�o�o�o�o �o�o�OV�O1 u����
��� ��)�;���_�q��� ������ˏݏ�<���%�r�I�[�m����$�DCSS_PST�AT ����ӑQ  �  �� � (�+��O���t� r�Ԑ�������������ӕ����կ�ĔSETU�P 	әB�������8�R�ͬs��b���������T1SOC 2
+������Cz������صCoP R�D�DLj�|�>�ϲ��� ���������0�B�T� #�xߊ�Yߛ����ߡ� ������>�P�b�1� ����y������� �(���L�^�p�?��� ��������������$ 6Zl~��Vϫ �D���); Mq��d�� ��//�7/I/[/ *//�/�/r/�/�/�/ �/?!?�/?W?i?8? �?�?�?�?�?�?�?�? O/OAOOeOwOFO�O �O�O��O�O_�O+_ =_O__s_�_�_f_�_ �_�_�_oo�_9oKo ]o,o�o�o�oto�o�o �o�o#�oGYk :������� ��1� ��g�y�H� �����������	��O -�?�Q�؏u�����h� ��ϟ������;� M�_�.�������v�˯ ݯ�����%���I�[� m�<���������ٿ� ��̿!�3��W�i�{� Jϟϱ��ϒ������ ��/�A�S�"�w߉�� j߿��ߠ������� =�O�a�0����x� �������'���K� ]�o�>����������� ������#5Yk }L������ �1Cgy� Z߯��Z�	// �?/Q/c/2/�/�/h/ z/�/�/�/??)?�/ M?_?q?@?�?�?�?�? �?�?�?O%O7OO[O mOONO�O�O�O�O�O �O�O�O3_E__i_{_ �_\_�_�_�_��_o o�_AoSoeo4o�o�o jo�o�o�o�o+ �oOasB��x �����'�9�� ]�o���P�����ɏ�� ���Ώ#�5�G��k� }���^���şן���� ���_C�U�ܟ6��� ��l���ӯ寴�	�� -���Q�c�u�D����� z�Ͽ��¿�)�;� 
�_�qσ�RϧϹψ� �������%�7�I�� m�ߑ�`ߵ����ߨ߀�����3�E�W�&���$DCSS_TC�PMAP  ������Q_ @ .�.�.�.���.��.�.�.�	.�
�.�.�.�.��.�/�  .��.�.�.�.�J.�.�.�.�.�U.�.�.�.�U.� .�!.�".�U#.�$.�%.�&.�U'.�(.�).�*.�U+.�,.�-.�..�U/.�0.�1.�2.�U3.�4.�5.�6.�U7.�8.�9.�:.�U;.�<.�=.�>.��?.�@u�UIROw 2��������������� ,>Pbt���@����-��� -��Qcu��� ����//)/;/ M/_/q/�/�/2�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O�/3O�/WOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_�&O�_q�UIZN �2��	 ��� �� oo$o*��_Rodo vo9o�o�o�o�o�o�o �o*<Nr� �Y������ &�8��\�n�=����� ��ȏ������ߏ4� F�X��|�����o�ğ ֟蟫���0���T� f�x�;�M�������������_x�UFRM� R�����8 1�^�p�/����ʿ ܿ�� ���6�H�#� l�~�YϢϴϏ����� ���� �2�I�V�h�� �ߞ�y����߯���
� ��.�@��d�v�Q�� �����������*� A�N�`������q��� ��������8J %n�[���� ��"9�FX� |�i����� /�0/B//f/x/S/ �/�/�/�/�/�/?? 1(?P?b?=?�?�?s? �?�?�?�?O�?(O:O O^OpOKO�O�O�O�O �O�O __)?;?H_Z_ �O~_�_k_�_�_�_�_ �_�_ o2ooVohoCo �o�oyo�o�o�o�o
 3_@R�ov�c �������*� �;�`�r�M������� ̏ޏ����+8�J� �n���[�������ǟ ���ٟ"�4��X�j� E�����{�į֯���� ��