��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ̊c��AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@ � �ALRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �� PCOU�PLE,   �$�!PPV1CESI0�!H1�!�PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q�!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W�1�W 6P�!SBN�_CF�!�0�$!J� ; 
2�1_�CMNT�$F�LAGS]�CH�E"$Nb_OP�T�2p�(CEL�LSETUP 7 `�0HO�0 �PRZ1%{cMAC{RO�bREPR�hD0D+t@��b{�e[HM MN�B
1^�UTOB U��0 9DoEVIC4STI�0��� P@13��`B�Qdf"VAL�#IS�P_UNI�#p_�DOv7IyFR_F�@K%D13�;A�c�C_WA?t�a�z�OFF_@N�DEL�xLF0q�A�q�r?q�p�C?�`�A�E�C#�s�A�TB�t�d�MO<� �sE � [�M�s��2�REV��BILF��1XI�� %�R  �� OD}`j�$NO`M�+��b�x�/�"u�� ������!X�@Dd� p E RD_�Eb��$FSS�B�&W`KBD_S�E2uAG� G�2B "_��B�� V�tp:5`ׁQC ��a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR�� BIGALLOW� (KD2�2�@VAR5�d!�A�B e`BL[@S �C ,KJqM�H`S�p�Z@M_O]z��w�CFd X�0�GR@��M�N�FLI���;@UI�RE�84�"� SW�IT=$/0_No`S��"CFd0M�{ �#PEED��@!�%`���p3`J3t	V�&$E�..p`|L��ELBOF�  �m��m�p/0��C	P�� F�B����1x��r@1J1E_y_T>!Բ�`��gt���G� �0WARNMxp�d�%`�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�M�� R�r$OR�I�.&ӧRT�S�Fg��CHG*V0I�p�T��PA
�I{�T�!��>� � �#@a����HDR�B��2B�BJ; �C��3�U4�5�6�7օ8�9>���x@�2w @� TRQ���$%f��ր����_�U������Oc <� ����Ȩ3�2^��LLECM�-�MULTIV4�"$���A
2q�CHILD�>�
1��z@T_1b � 4� STY 2�b4�=@�)24�p���@�� |9$��T�A�I`�E���eTO���E��EXT���ᗑ�B��2G2�0>��@���1b.'��B ��A�K�  �"K�/% �a��R���?s��=�O�A!M��;A�֗�M�� 	�  =�I�" L�0[�� R�z�pA��$JOBB������`���IGI�# dӀ����R�-'`r��A�ҧ��_M�n�b$ tӀFL6��BNG�A��TBA � ϑ�!��
/1�À �0���R0�P/p ,����%�|���Bq@W�
2JW�_RH�CZJZ�_zJ?�D/5C�	�ӧ���@����Rd&A������ȯ�qGӨ�g@NHANC��$LG/��a2qӐ� ـ�@��A�p� ���aR���>$x��?#DB��?#RA�c?#AZ�t@�(.�����`FCT����_F࠳`�SM��!I�+lA�% ` �` ���$/�/�@���[�a��M�0�\��`��أHK��A�Es@͐�!�"W��Nz� SbXYZW�`D�"����6��C�����'  . I�I��2�(p�STD�_C�t�1Q��US�TڒU�)#�0U�[�%?IO1��� _Up�q�* \��=�#AORzs8Bp�;�]��`O6  RSY�G�0�q^EUp��H`�G�� ��]�DBPX�WORK�+���$SKP_�p��D�B�TR�p , �=�`����Z m�bOD3��a _C"�0;b�C� �GPL:c�a��tőS�D�W��3Bb����P��P M)DB�!�-�B APR��
�@Ja3��. /�u����� �LuY/�_�S���0�_���PCr�1�_�TENEG��]� 2�_�SVPR�E.��R3H {$C��.$L8c�/$uSނz IkIN�E�WA_D1%�ROyp�������q�c�7 t@�fPA���R�ETURN�b�M�MR"U��I�CR�g`EWM@�SIGNZ�A ���e�� 0$P'�g1$P� m�2pB�p'tm�+pD�@� �'�bdNa)r�GO_AW ��@ؑ�B1�@CSd�(�C%YI�4���`1w�qTu��t2�z2�vN��}��E}sDEVI�s` 5 P M$��RB��I�wyPk��I_BY����"�T7Q�tHND=G�Q6 H4��1��w��$DSBL C��o��vg@�Ʈ@qL��7O�f@]���3FB���FEra8��ׂ�t}s���8> pi�T1?���MCS����fD �ւ[2H� W ��EE���%F����t����9 T�p��x�NK_N:�����UZ��L�wHA�vZ' ~�2���P~r�q7w: �=MDLn���9�ጂٱh����! e����J��~� +����,�N�D����3���ՒG!aqSL�Ad�7;  ��INP��"�����}q_ V�4<�06`C� �NU��  D�L�ק��SH!�7=BM��q���ܢӢ����g���>P +$ٰ�٢��^��^�Y�FI B�\��Ă��'A	'AW�l�NTV��]�V\~�X�SKI�#T� ��a�ۺ�T1J�3:39_�P�SAFN����_SV�EXCSLU��N@�DV@�Ll @�Y����S�H�I_V
0\2PPL5YPRo�HIM�T��n�_MLX��pVORFY_�Cl�M��gIOC�UC_� �����O�q�LS(�0v�FT4Q���)��@P�E$�t��A��CNFt�6եup��pm�4ACHD��o������AFC C	PlV�TQTP?�� ί� ?`�@TA��@�0L@ ��N���]� @����T��T! S����te@{R�A DO�� w23���!n��	_1�#�H!�̔�΀�K��B�2��MAR�GI�$����A ���_SGNE�C;
$�`�a^aR0 ��3��@ B��B��ANNUN�P?����uCN@�`%0��`��� ���BEFc@]I�RD @Q�F���4OT�`�sFTӠHR,Q��CQ0�M��N�I|RE�����A�W���DAY=CLOCAD�t;T|�<S5}�EFF_AXI��%F`1QO3O��Eq���@_RTRQ�E�G����0RQ
j�Evp ��|��F�0f�R0 �tp��AMP�E<� H 0�`œ^��`Ds�DU�`��v�BCAr� I?��`N ErIDLE_PWRI\V!n0�V�wV_[ |�� ��DIAG�5J�o 1$V�`SE�3TQl�e��P�l�^E_��j�VE6� �0SWH�q (� �b|�Gn�3OHxPPHk�IRAl�B�@�[� �a�bk��w3�O  � ��v�|�I�0 ��pRQDW�MS-�%AX{6j�LIFE�@�&�MQy�NH!Q%��F#�C����CB0�mpNr$�Y @�aFLAl�f��OV0]&HE��>l�SUPPO�@u��y��@_�$��!_�X83�$gq�'Z�*W��*B1�'T�#`�k2XYZáj�Y2D8CY`T@�`N�����f� �C�k���IC�TA�K `�pCACH�ӫ�3�����I��bNӰUFFI� \��@��;T��r<S6CQ.�MSW�5�L 8	�KEYI7MAG�cTMLa���*Ax�&E���B��OC�VIER-aM ���BGL����y�?G� 	��П4N�m:�ST�!�B P�D,P�D��D��@�EMAI䐔a��p��r�FAUL|RO bB�c�� spUʰMA�"`T'`E�P< �$S�S[ � ITw�BUF�7y��7r�tN[�LSUB1T��Cx�o�R�tRSAV|U>R'c2�\�WT���P�T�*`S�n�_1PbU���YOT(�bK��P��M��d����WAX��2��X�1P��S_GH#
$��DYN_���Q� <Q�D��0����M�� T�F��`|�\�DI��EGDT_Pɰ:�R��b�GRQM�&��Jq�a����׀��Fs� 7S (�SVqpB���4�_�.��a��T� �@���B�S7C_R]1IK>B'r��$t��R"A#u�H�a'DSP:FrP�lyIM|Sas�qz��a� �U>w� <1%sM�@I�P��s��0`tTH�b0ЃTr��T`asH9S�cCsBSCʴq0�� V�����S�_�D��CONVE�G ���b0^v1PFHy�adCs�`&a?ASC����sMERg��aF�BCMPg��`ETn[� UBFU� DU%P�D�:12��CDWy�p�P�CG�&[@NO6�:�V� �H�� ���P���C�����w��A��`���WH *�L Ơ�Cc�W����Y�� ���р�q�|��񨀖A��7}�8}�9P}�H ���1��1��U1��1��1ʚ1ךU1�1�2��2�����2��2��2��2�ʚ2ך2�2�3J��3��3����3��U3��3ʚ3ך3��3�4��QEXT[�X[b�H``t&``�z�k`˷$���FD�R�YTPV���RK"	��K"RE�M*F��]"OVM�:s/�A8�TROVf8�DT�PX�MXg��IN8ɉ W��IN	Dv�["
�ȕ`K ^`�G1a�a��@Q%7Da�RIV��u"]"oGEAR:qIO.	K(�[$N�`���,(��F@� \#Z_MC�M<0K! �F� U�T���Z ,�TQ?' b�y@t�G?t�E |�.�>Q����[ �Pa� RI�E���UP2_ \ ��@=STD	p<TT����������a>RBACUb] T��>R�d�)�j%C�E��0��IFI��0��i�{�4��PTT��FLUI�D^ �?0gHPUR�gQ�"�r�a��4P+ I�$��S�d�?x��J�`C9O�P�SVRT��N�x$SHO* ��CASS��Qw%�pٴBG_%��3�����FORCx�B��o�DATA��-_�BFU_�1�bb��2�en�b0��` |�K`NAV	`�������$�S�Bu#�$VISI���2S�C	dSE�����VZ��O�$&�BK�x�� ��$PO���I��FMR}2��a � �	��`#��&ߠ8�O� (�_����+IT_^�ۄ)�M�����DGCL�F�DGDY�L	D����5Y&��Q$YѩM됇CbN@{	� T�FS�P�Dc� P��W�cK $GEX_WnW1%`�]��"X3�5��9G+�d �K`���SWeUO�DEBcUG��-�GR�к;@U�BKU��O�1R� _ PO@_ )�����M��gLOOc>!SM� �E�R�a��u _E �e >@�G��TERM`%fi'O�ORI�ae gi&��`SM_�`>Re h�i%V�(ii%3U}P\Bj� -��F�e��w#� f��yG�*ELTO�A9�bF�FIG�2�a�_���@�$�$g$U;FR�b$�1�R0օ� OT_7F�TqA�p q3NST�`�PAT�q�0�2PT�HJ�ԀE�@�c3ART�P'5�Q��B�aREL�:�aS�HFT�r�a�1�8_���R��у�& � $�'@i�
����s@b�SHI�0�Uy� �QAYLO�p�Oa�q�����1����pERV��XA��H��m7��`�2%�P�E3�P�RyC���ASYM�a���aWJ07����E �ӷ1�I��ׁUT�` Oa�5�F�5P�su@�J�7FOR�`M  �O!k]��5&0�0L0���HOL ;�l �s2T����O�C1!E�$�OP��qn���H$�����$��PR^�f�aOU��3e���R�5e�X�1 �e$7PWR��IMe�BR_�S�4�� �3�aCUD���`�Q�dm���$H�e!�`AD+DR˶HR!G�2�a��a�a ��R��[�n H��S����%��e`3��e���e��SEl��L�HS�MNu�o���Pªq��0OL�s߰`ڵ�I ACRO��&1��ND_C�s��Afd�K�ROUP��R_�В� �Q1|�=�s ���y%��y-��x���y���y>�=A��Ҁ�AVED�w-��u�`<(qp $���P�_D�� ��'rPR�M_��HTT�P_�H[�q (�ÀOBJ��b �$˶LE~3�P��\�r � ���ྰ%_��TE#ԂS�PIC��KRLPiHITGCOU�!��L�� �PԂ������PR��P�SSB�{�JQUE?RY_FLAvs�@_WEBSOC��G�HW�#1��s�`}<PINCPU(���O���g�����d�t��O��IO�LN�t 8��R���$SL!$INPUT_U!$`��Pw�֐SSL.���u����2�.��C��B�IO^a�F_AS=v��$L+ਇ+�A ��bb41�����Z@�HYʷ����#qe�U;OP:w `v�ϡ�˶�¡�������"`P IC`���� �	�H��IP_ME��v�x Xv�IP�`(�R�C_N�p�d���R0ʳp�ױQrSP �z��C��BG(� ��M��Av�y lv@CTiApB��AL TI�`3UfP_ ۵�0PSڶBU_ ID� 
�L �� `�a�����0�z)����ϴ�N�N�_ O��IRCA�_CNf� { ��Ɖ-�CYpEA��������IC����tpR�=QDAYy_
��NTVA������!��5����SCAj@��CL�
����
���v�|5�VĬ2,b�l�N_�PCV�n�
���w�})�T��S�р���
��e���T� 2| $� �v��~��֣�ذLABp1��_ ��UNIX�9�ӑ ITY裪��e��p�� ��<�)���R_URLn���$A;qEN ����s`vsTeqT_�U���J��X�M�$���E�ᒐR�祪�� A�,���J�H���FLy��= 
|���
�UJR|U� ���F�6G���K7��D>�$J7,�s��J8*�7���$3�E�7��&�8\�)�oAPHIQ4�zy�DkJ7J8Rޒ�L_KE'� o �K͐LMX�� � <U�XR�i�����WATCH�_VAZqu@AំF'IEL`��cyn���&:� � u1VbwP�CTX�j�����LGE���� !��LG_SIZ΄�[8Zm�ZFDeIYp1! gXb ZW �S`� 8�m��� �b ���A�0_i0_CM c3#�*'FQ1�KW d(V(Bbpo pm�p� |Io�1 pb p�W RS��0  M(C�LN�R�۠-�DE6E3��� �c�i���PL#�7DAU"%EAq�͐�T8". GH�R��y��BOO�a��3 C��F�ITV�l$�A0��RE���(SCRX����D&�ǒ�qMARGI4�Sp�,@����T�"�y�S���x�W�$y�$��JG=M7MNCHt�y�FN��6K@7r�>9�UFL87@L8FWDvL8HL�9STPL:�VL8"�L8s L8RS"�9HOPh;��C9D�3 R��}P�'IUh�`4@�'�5$ ��S2G09�pPOWG�:�%�3,�64��N9EX��TUI>5I� �ӌ���� �C3�C<0'�,�o�:��&�@�!NaqvcAcNAy��Q�AI]�8gt7Ӝ�DCS���c�RS�cRROXXOdWS��ÂRoXS{X�(IGNp 
Ђ=10 ��[T�DEV�7LL���; B��C �	 8�Tr$f/蛒����Z�3A�a�	 W�h萦�Oqs�S1Je2Je3Ja��BSPC G� �ƋG`-T� �%��Q�T�r@�&E�V�fST�R9 YBr~�a �$E�fC�k�g��f	v9�CB� L����� �� u�xs뀔�g�q�jt���!�#_ ����ʐv�#Ӡ �s �M�C�� ���C�LDP᠜�TRQ�LI ���y�tFL ���rQ��s5�D���w�~�LD�u�t�uOR�G���1�RESERV��M���M�Œ��t��� � 	0�u�5�t�uSV��p���	1�����RCLMC��M�_�ωА���_C�MDBG�h�I����$DE?BUGMAS�������U�$T8P��EtF�d��pFRQҤ�� � K	H_RS_RU4�bq��A��$EFREQ�6u!$0YOV�ER�k��f�PnU1EFI�%GqȤ� �
Y�z�� q\����E�$U�`Ρ�?��
�PSI`��	��CA ��ʲ��σUY�%�?({ 	��MISC��g� d��aRQ���	��TB� � ���A��AX���>��EXCESg�9Rd�M�H�9�u�؜�}qd�SC�` '� H�х�_������������pKE䔰�+�� &�B_, F�LICBtB� QU�IRE CMOt�O���얩qLdpMD� �p{!��5b���$L�MND!���I����L �D|;
$INAUT�!�
$RSM�ȧPN��b�C���PS�TLH� 4U�L�OC�fRI"��eEX��ANG.R.����ODA]��q��� �RMF0�����icr�@mu���$�S�UPiu��FX��I�GG! � � ��cs�F�cs
Fct�� ޒ�b5��`E��`T�5�0tC��g�TI��C`�;��M���� t&�MD���)��XP���ԁ��H��.���D#IAa��Ӻ�W�!�Ԩ0af���D@#)֡O��㥀��� �C�Up V	���.���Or�!_��� �{`0�c������ |�P|��0� ��P{�KqEB��e-$B��o�=pND2ւ�����2_TXltXTR�AXS������LO�: ����}�L����C�.�&�[�R�R2h��� -��!A�� d$OCALI���GFQ:j�2F`RINbn�w<$Rx�SW0ۄܨ��ABC��D_�J��{�q��_J3:��
��1SP, �q�P����3��H�9p
q�#J�3n����O�QIM耯�CS�KP�zb7?SbJ+ᯂQb�y�����_AZ��/�E�L�Q.ցOCMP0�ð�� RTE��� �1�0 ���1���@ ZSMG��0�Э�JG�pSCyLʠ��SPH_�P���f��q�u�R'TER��n�Pk�)_EP�q�`A� �c̯��DI�Q23=UdDF  ����LW�VEL�qIqNxr�@�_BLXP.��Y/�J��'>$  �IN���B]�C�9%�".�8!:6p_T� �F%a"���^$��k)�~p�DHʠ��\�9`�$Vw��_�A$�=��~�&A$���S�h��H ��$BEL� m��_oACCE� 	8<�0IRC_�q��@�NT��c$SPSʠ�rL��� M4�s9 .7��GP/6��9�7$3�73S2T�͡_Ga�"�0�1��8�17_MG}�DD�1�~�FW�p��3�5$3�2�8DEKPPA�BN[7ROgEE �2KaBO�p�Ka���1�$USE_tv�SP��CTRT�Y4@� �� <qYN�g�A�@�FR �ѢAM:�N�=R�0O�v1�DINC(��B�4����GY��ENC�L���.�K12��H0IN¿bIS28U��ONT|�%NT23_�~�fSLO�~�|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1����PERCH  �S��� �W���SlщR ��l����E�0�0P	AS2EeL�DP7�O�NUЉZ�f�VTRK�RqAY"�?c��a S2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gBT��DUX �2S_BC?KLSH_CS2Fu :��V���C-�esRoz|�A�CLALMJTp@��`� �uCHKe |����GLRTYp� ��8T��5���_�ùT'_UM3��vC3��1�Z���LMT��_ALG��%���0�E*� K�=�)�@5F�@8 9��Nb��)hPC�Q)hHpТ��5�uCMC��\�0�7CN_��N��L�;SF�!iV�B���.W���S2/�ĈCAT�~SH�Å��4  V�q/q/V�T1�f�0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e��R� @B�_Wu�d@�!a��#`��#`�Ih�Iv�I�#F��S�:X��I�0VC00��֢1ܮ�0�⦇JRKܬ!��<�D�BXMt�<�M�_sDL�!_bGRVg�``��#`��#A�H_%�8?��0��COS��� ��LN#���ߥŴ�  ��=������꼰�<�1Z���VA�MYǱ:���᯻[�THET=0�UNK23�#��l�#ȰCB��CB�#Cz�AS�ѯ����#����SB�#��'GTSkZAC�����&���$DU�phg6�j��E�%eQ%a_��x�NEhs1K�t�� y��A}Ŧկ׍�����LCPH����^U��Sߥ ����������!��(Ʀ�V��V�غ ��UV��V��V
�V�UV&�V4�VB�H��@������d�����H
�UH�H&�H4�HB�O��O��Os���O���O��O
�O�O*&�O4�O(�F�Ҫ��	���SPBA?LANCE_J�6�LE��H_}�SP�>!۶^�^��PFULCb�q����K*1�UTO_<�p�uT1T2�	
22N�q2VP�M�a�� i�Z23	qTu`O��1Q�INSEG2�QREV�PGQgDIF�ep)1�U6�1��`OBK�q�j�w2,�VP�qI�L�CHWAR4B�BA�B��u$MEC�H��J��A��vAX��aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ�@��C1_ɒT �� x $WEgIGH�@�`$��d\#��I�A�PIFvAN�0LAG�B��S�B�:�BBIL�%OD��`�Ps"ST0s"P:�pt � N�C!L ��P 
P2�Aɑ � 2��Tx&DEB�U�#L|0�"5�M'MY9C59N��$4Ώ`$D|1 a$�0ېl� > D�O_:0AK!� <@_ �&� �q�A��B�"�� NJS�8_�P�@���"O�p ��� %�T7P?Q�TxL4F0TICK�#�T1N0%�3=p�0!N�P� u3�PR\p�A��5��5U0PRO�MP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a�@�RU�COD�#FU�@�&ID_�P�E8�2B> G_SUFF��� �#�AXA�2DO�7/�5� �6GR�#��DC�D���E��E-��DU4� ��_ H_FI�!�9GSORD�! R 236s�HR�AN0�$ZDT�Et�p�!X5�4 *WL_NA�1�0�R>�5DEF_I�X�R F�T�5�"�6�$�6�S�5�UFISm�#�m1|��40c�3�T6�44􁆂�"D� ?rfd��#D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D �S�D�U�D>b�B�c�E �S�Dd�B�&2v2a�C �ʑ�E�R�E�S�C9wwu�H�0P} d�0,aĂ�F0W�h�u�c4�80�TE�qY4�� �!LOM�B_�r�w0s"VI]S��ITYs"Aۑ}O�#A_FRI���~SI,a�n�R��07��07�3�#s"WB�W�Q��%�_���AEAS{#�B��P|�x`WB8�45�55��6|#ORMULA�_I���G�W�� h 
>75C?OEFF_O�1&H)��1��Go�{#S� �52CA� :?L3�!G�Rm� � � �$�`�v2X�0TM�g���e�2�c��3�ERIT�d�T� ��  �LL�Dp`SΛ�_SVkd��$��v� �.���� � ���SETU,cMEAG@�@Πt �!HR>L � � (�  0��l��l��aDw��R�0�a�a}d�]�d��B��Ay`�Gax`��[Ѐk@R�EC[Qq�R0MS�K_A y�� P~_!1_USER������*���VE�L����-�!��I�zPB�MT�1CF}G���  �0z]O�NOREJ �0l���[�� �4 e���"�X�YZ<SB� 3�0ށ�_ERRK!� U ѐ�1�@c�Ȱ�!��>�B0BUFI�NDX��R0� MO�Ry�� H_ CU ȱ�1��dAyQ?�I�>Q$ +��a����� \�G{�� � $SI�0h��@2	�VOv�qО- OBJE| w�A�DJUF2yĈ�AYh�����D��OUKPp����AMR=��T��-���X2DI�R����Xf�1  D#YNt�0�-�T� ���R��0� ���OP�WOR�� �},B0SYSBU����SOPo���zډUy�XP�`K���P�A�q������OP
�@U���}�"1^��IMAG۱_ ��п"IM.���IN�������RGOVR!D"ё�	���P����@  >gplcC��L�`�BŰ?l�PMC_QE�P�1N��Mr��1212R�"�SL�| ��� �R OV�SL=S�rDEX�\a`��2�:�_ "���P#���P������2�C �P>���#�_ZERl�8��:���� @��:��O�@RIy��
�[�g@e���s�P�PL����  $FWREEY�EU�~�TZ��L����T��� ATUSk�,1C#_T�����B�������p�Vc1��P���C Dc1�к���LQ�����MQ��ۡL�XE@��x�5IP�W��` ��UP��H`&aP!X;@��43�����PGY��g�$SUB���q�����JMPWAIT8~ ���LOW���1wē CVF_A�0�b�R�Z��CC ��R$��28IGNR�_PL��DBTB2� P*a�BW@.2t�U�0-IG��!@=I�TNLN,��RBѡb�N!@��P�EED~ ��HADCOW� ��t���E��p����PSPD��� L_ A�нP���	#UNq � �RP (�LYwPa��}��PH_PK����b�RETRIE���x���2�R!D@FI��� ���V �$� 2�d�DBG�LV<LOGSIYZz�baKTU��r�$D��_TXV�EM�Cڡ)�� �-�R�#�r��CHECAKz����L���ϰ�q)�L��NP�A�`TJ"����)1P4����
�AR�"�BC =Sa��O�@����ATTS�u䡳&� 0w�^a�3-#UX^�4��PL�@Z�� $�d��qSWITCH��h�W��AS���f�3LLB���� $BA�Dvc��BAMi��6I��(@J5��N�UB�6[F
A_KNOWhK3qB"�U��AD+H�c� D��IPAYGLOAq�9p�C_����GrѼGZ�CLqA�j��PLCL_6� !4��BOA?�T*7�VFYCӐ�J(p��D�I�HRՐ�G$�TB��6�J(�zQ�_J�A �B�AN�D����T�BQ������PL@AL_ ��0 =�TATe��pC��D�CE����J3�P�V� T�PDCK^�)b���COM�_ALPH�ScBE<�߁�_�\��X�x\� �s ���OD_1�J52�DDM�AR<�h��e�f�cQ�TIA4�i5�i6��MOM�(��c�c�c�c�cV�B� AD�cv�cv�cPUBP�R�d<u�c�<u�b}"�1���� L$PI$��pc@��G�y��I�yI�{I�{I�s�`�A���v��v�J�b��a��HIG�3�� �0���5�0�f��?�5N�5�SAMPD Ƣ�0����;@�S ��с6��� 1���� ���`���`�1�K�P��`腽P�H��IN1��P��8� T�/��:�z�Q�z���/GAMM&�S��$GET������D^d>�
$�PIB�R��I��$HIB��_���1��E=�b�A�9�*�LW� W�N�9�{�*�Zb��:�QCdCHK0�j�ݠnI_��M�J� �Roh�Q ��sJ�-v|��S �$�X� 1�N�I�R�CH_D$R1N���^�LE���i�p�Zh8�ţMS�WFL/M�PSC�R�75�Ҽ ��3 �"Ķ�6��`��ع��紙��0SV���P'������GRO<�g�S_SA=AH�,=ńNO^`Ci� _d=��no�O�O�x������p�B�u�ȐcDO�A��!�ں�*� t�:�Z1f�;�7����C� �Q�0Mmu� 7� �YL�snQ ��� ���"��<s�	�����nQ૰�<3M_Wl��� ��\p��(�o�MC��P���Q�����hpM.�pr� ���!��$�WM��ANGL�!�AM�6dK�=dK�DdK��TT7�N�k@��3�#�PXC O�Ec�QZ��hp	nt�[ ���OM��� ϑϣϵ����`� c��Z0j�^a_�2� | a�J��i���c���c�J��j�����jA� P���{���  �@�{�P�1�PMON�_QU�� � =860QCOU��7QTHxHO��B 7HYS�0ESPBB �UE- 3�f0O�4΋  c P�^�R�UN_TO�� 8o ��� P�@�<�INDE�#_PGGRA���0��2�ПNE_NO��I�Tf��o INFOB��a"�����P!�OI� (*�SLEQ!�*�*��&S��l4� 4�60ENABy� PTION�3��r���^GCF�!� �@60J�Q���R�d!��
�P�EDIT�� ��� ��KAQ"� �E�(�NU'(AUT<Y�%COPYAQ�(2,�qe�M�N< @+^��PRUTm� C"�N�OU�2$G���$#RGADJZ��u2X_��IX�P���&���&W�(P�(�~��&9�� 
�N�P_�CYCy�H�RG�NSc�{�s�LG�O£�NYQ_FREQSrW@��X1�4�L�@�2P0�!�c@�"�CRE��Mà�IF�q�NA���%�4_Gf�STA�TU~�f��MAI�L��|CIq�=LA�ST�1a*4ELE�Mg� ��QrFEASIt;�ւΰ ��B"�F�AF����I� ��O2�E u�&vBAB��PE� =��VA�FzQ�I��TqU�[��R��S�FRMS_TRpC�Qc� �C��Z�
��1�D�*4�ns؆�	MB 2� `���N�3V �R2WR*���шR^W��wj�DOU�^�NL�,2PR`�h�1�GRID��BARS!�TYuZ��Op�� |_"�4!� �R�TO��d�� � ����P�OR�c~vbSReV�0)"dfDI[�T�`;aNd�pXg
�XgQ4Vi��Xg6Vi7ViI8:a�Fʒg�z ?$VALU�C0��3D�� F05��C !pT���S�1�-ȆAN/��b�1R��]11ATOTALX����=sPWE3I�Q>StREGENQzfr��X�H�]5	v( cTR�CS�Qq_S3��wfp�V�!��r��BE�3�PG0B�( nsV_H�PDA(��p�S_Ya���i6�S��AR(�2� }�"IG_SE�3ȿpb�5_� �tC_��V$CMPl��D�Ep�G���IšZ�~�X��R�aENHA{NC.� p Q�r�2���INT�9`cq�F���MAsSK�3�@OVRMP �PD�1-��W��c�U�l�_RF�{�V��PSLGP�g��9�j5��,�;pDpqS���4��U�������TE���`�#��`k���J^�Y�y3IL_Mx4�s��p��TQ( ���@ԍ���V.�C<�P_h �R�F�M]�V1\��V1j�2y�2j�3*y�3j�4y�4j����p۲������ܲIN�VIB8�6�#�T�*�2&�22�3&�32�4&�42��6��|�J�  �T �$MC_FK `�� �L>�J�х1pMbj�Iу��zS ���1���KEEP__HNADD��!�$�@�C��0	��Q����
�O!�v ��p�p
�և
�REM!	�Cq�RF�]�b�U��4e	�HPWD w �SBM��~�PCOLLAB*��p��/q�2IT�/0��Q"NO1�FC�ALp⎵��� ,� �FLv�A$SSYN���M��Ck���RpUP_DLYz��zDELA9дDq�2Y AD(����QSKIPO��� �`� O��NT����c�P_� ��� � ��cp���q�ٞ�� o`��|`�ډ`�ږ`��У`�ڰ`��9�!�JS2R0  �lX�@TR3H��1AH� �pH����`RDCq���� � R�R, 5��R�1��E��5TRGE�_C��RGFLG"���W��5TSPC�1UM�_H��2TH2N�}Q�;� 1� �;��Q02 � D� ˈ��@O2_PC3W�S��|�1Y0L10_Cw2q��,��� � $\� U@��V7�@����0��VU \����� rd��C� �+��7��DZ G\s�RUVL1[�1h����10]�_DS`�������PK 11�� lڰ����q��AT?��$�Q[7� � ��K 5T���oHOME� ��
c2h�n���(���3h���0!3E *�c4h�hz���(�&0`5h����	//-/?/Q'6h��b/t/�/�/�/�/�7h��/�/??'?9?S ���!8h�\?`n?�?�?�?�? _�S����  p�Aa{p����+�z_�Ed� T=�nD4vnCIO䑎IIt@`�O��_OP�E�C.r���POWE	�� X@�f� �$$Cd��S����j@���3�3� �@�S�I��GP�0�QIRTUA�L�O
QAAVM_�WRK 2 7U� 0  �5Qn_zX�k_�] �\	 �P�]�_3�8P��_�_�Ve�\#m/o�Q5o0jo|o�dHPBS��� 1Y� <Xo�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ�b�C$�AXLM�@v���c  d��IN����PRE�
�E�J�-�_U�P��[�7QHPIO�CNV_�� �	�Pr�US>��g�c{IO)�V 1U[P $E`��Qս9lҿ8P?�� ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o��o�m�LARMRECOV a���-���LMDG ���ɰ�LM?_IF ��� ை����zv����%�6�, 
 6�_��r漅�������̍$w���׏���8�J�\�n����NGTOL  a�� 	 A   ���ț�PPINFoO ={ <v�����1��   I�3�a�"rP���t��� �����ί���>�o����j�|������� Ŀֿ�����0�B��PzPPLICAT�ION ?����+��Handling�Tool �� �
V9.30P/�04ǐM�
88g340�å�F0����202�ťʚϬ�7DF3��M̎��NoneM�F{RAM� 6���Z�_ACTIVE��b  sï�  ~p�UTOMODz��A���m�CHGAoPONL�� ���OUPLED 1ey� �������g�CUREQ �1	e{  T�
��	p��w����#r���e�HN���{�HTTHKY��
$r��\[�m���� O�	�'�-�?�Q�c�u� ������������ #);M_q�� ����% 7I[m��� /���/!/3/E/ W/i/{/�/�/�/?�/ �/�/??/?A?S?e? w?�?�?�?O�?�?�? OO+O=OOOaOsO�O �O�O_�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_oo#o5o GoYoko}o�o�o�o�o �o�o1CU gy������ �	��-�?�Q�c���1�TO��|�p�DO_CLEAN��|n��NM  �� �B�T�f�x����%�DSPDRY�R��m�HI���@ /�����,�>�P�b��t���������ίj�MAXa�ۄ��������Xۄ������p�PL�UGG��܇�ӌ�P�RC��B� ���ׯF�OK���ȔSEGF��K������ �.�����,�>�v���LAPӟ澨�� �϶����������"��4�F�X�j߯�TOT�AL�7���USE+NUӰ�� �������1�RGDISPWMMC����C��&��@@Ȓ��Oѐ������_STRI�NG 1
��
��M��Sl��
A�_ITEM1K�  nl�g�y�� �����������	�� -�?�Q�c�u����������I/O S�IGNALE��Tryout M�odeL�Inp���Simulat{edP�OutOVERRА� = 100O�In cycl�P�Prog A�borP���S�tatusN�	H�eartbeat�J�MH Fauyl��Aler�	 ������*8<N` ׃G� ׁY�c����� ////A/S/e/w/�/��/�/�/�/�/�/wWOR��G�-1�?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO8�O�O�NPOE� �@E;�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo�BDEV�Nu`�Obo�o �o�o�o�o�o, >Pbt��������PALT ��E?�A�S�e�w� ��������я���� �+�=�O�a�s����GRI�G뽑1��� ���	��-�?�Q�c� u���������ϯ�� ��)�����R�a� ՟;���������ѿ� ����+�=�O�a�s���ϗϩϻ���O�PREG��y���-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_��q����$ARG_�-0D ?	������� � 	$��	+[��]����������SBN_CONGFIG���� ��CII_S?AVE  ��)����TCELLSETUP ���%  OME_I�O����%MOV�_Hn�����REP�d�����UTOBA�CKY���#��FRA:\�� �����)�'`l ���&� 7"�� 24/0�6{  09:35:24�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� ,,		�����O�G�O __#_%_7_q_[_�_ _�_�_�_�_�_�_%o����D�@TSK � �M&,O��UP3DT�@EGd�`�F�XWZD_ENB8ED��fSTADE��ܖe��XIS�UNOT 2��&�(��� 	 0|�} Z�0&�? �<_ �/� K��pp�T<�bp�p�8t�}V��)q{|��t�� B=|�o���;9Յ�!{D�x�Q\��gMETc�2Lf�E� P qA|h�iA��A��B-��B��B�y��}?y�J�?��?:��&@5�W?U��s@���}S�CRDCFG 1��� ��z�����ԏ�����Q=���H�Z� l�~�����	�Ɵ-�� ��� �2�D���域���GR�`�`�O���0kNA����	��n��_EDC@1n��� 
 �%-�0EDT-q����L%�p��"���-������������^��  ����2����*�RIE���*� q���ϧ���3bϮ� @Ͻϯd?�����=�O���sϏ�4.ߞ�{��� ��W���	�߱�?ߏ�5��j�G����#�� ����}�6��6� �Z�����Z����I��7�����&��΀��&m������8^ҿ�����͇� 9K�o��9*�w����S��;��CR����B/ T//�/��w//���РNO_DEL�����GE_UNU�SE���IGAL�LOW 1���2p(*SYS�TEM*�s	$SERV_GR�;�B0�@REGK5$8m3�|B0NUMp:�3��=PMU� �u�LAY�p�|?PMPALD@�5�CYC10�.�>x�0�>CULSU�?0�=�2�AM3LOWD�BOXORIt5C�UR_D@�=PM�CNV�6D@1�0�>�@T4DLI��`=O_9	*PRO�GRAJ4PG�_MI�>�OPAL(�E_UPB7_B>�$FLUI_RESU�7p_z?�_�T#MRY>h0�,�/�b �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� ��������"�LAL_OUT �1;l���WD_�ABOR�0?d�I�TR_RTN  �����g�NONgSTOǠ�� 8�CE_RIA_IL0��ۀ��ŀFCFG ��x۔��_LIMY2�2ګ �  �� 	i�J��<�e�g��5��  9��������
����u��PAQPGP ;1�����Q�c�u�4�CK0����+C1��9��@���P�C��CV��]��d
��l��s���0����C[٤m��v���������� C�j���-���?�Â{HE� ONFI�P�q�G�G_P�@1� �%��������ǿٿ����G�KoPAUSaA1�ۃ �B�W��E� ��iϓϹϟ������� ���#�I�/�m��e�����M��NFO �1"��� �7��ߖ��C 	�=���?���h���'¶��ࠐ ��?��C�8��D�w�3�������B� h3�E�ŀO����c�COLLECT_�"�[�����EN�@��y���k�N[DE��"�3��"1234567890��\1��H ��֕H&��)M� r�\,L�^���]+���� ��������C 2 �Vhz���� ��
c.@R �v���������� ����I�O !���q����u/�/�/�/C'TR��2"'-(׀^)
��.R�#R-�*W�^ 9_MOR�$� �;�l5��l9�?r?��?�?�?�;E2��%JS=,W�?@�@��CR׀K)DցC�R��&u�XOWAWBC4 W A�q��׀x׀�A"@Cz  Bʇ@CG�B8��AC�  @yB�׀�ց:d�43 <#�
�E���I�OT�C=AI��'GM?�C��(S=���Qd=AT�_DEFPROG �;%�/m_APINUSE�V�ۅ��TKEY_TBL�  s�ہ���	
��� !"�#$%&'()*�+,-./�:;�<=>?@ABC�DPGHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����Ga���͓��������������������������������������������������?������!�P�LCK�\���P�PS�TAn��T_AUT/O_DO��NFs�IND���n��R_3T1wT2N�����5ŀTRLCPL�ETE���z_S�CREEN ~�kcscÂ�U��MMENU ;1)O� <�[_ #�q��,�a���>�d� ��t���ӏ����	��� ��Q�(�:���^�p� ������̟�ܟ�;� �$�q�H�Z������� ���Ưد%����4� m�D�V���z���ٿ�� ¿�!���
�W�.�@� ��d�vϜ��ϬϾ�� ����A��*�P߉�`� r߿ߖߨ�������� =��&�s�J�\��� ���������'�,�p_MANUAL��EqDB
12�v�iDBG_ERRLIPs*�{h! 0�������g�NUMLIM�s:QOE�@�DBPXWORK 1+�{��>P�bt��-DBTB_�q ,��kC3!�VD!DB_A�WAYo�h!GC�P OB=��A�_CAL���o�k�Y�p�uO@`�_�� 1-
�+@
-k-6[l��_M+pIS�`��@"@�ONTImM�w�OD���&
�U;MOTN�END�_:REC�ORD 13�{� ��[CG�O� f!T/[K��/�/�/�/ _(�/�/f/?�/??Q? c?�/?�??�?,?�? �?OO�?;O�?_O�? �O�O�O�O(O�OLO_ pO%_7_I_[_�O_�O �__�_�_�_�_l_!o �_,o�_io{o�o�oo �o2o�oVo/A �oeP^�
�� �R���=��a� s��������*�ߏN� ��'���ԏ]�̏�� ������ɟ۟v���n� #���G�Y�k�}����TOLERENC��B�0� L���g�CSS_CNS�TCY 24	�t���.����� �0�>�P�b�x����� ����ο����(��:�äDEVICEw 25ӫ � �ϟϱ������������/�AߟģHND�GD 6ӫ� C�zT�.!ơLS 27t�S������������/�U�ŢPARAM 8Gb��A�Ք�RBT 2]:8�<����CkA� �·�  � �A���.SB����A�B�  ����������.�����  ����A�A�C����c�u����C�A�D���k�pz�A�A��HA�c��A�	�?( uL^p���A��Bt/�D��C���_ 	 A�=��ABffA�#33AҊ��g�A�A�Cf���a��A�J��7B�]��B��B�ffBᴠ�3�3C$.@R� (����A��� �
/��//)/;/ �/_/q/�/�/�/�/�/ �/�/<??%?r?I?[? m??�?�?�?�?�?&O 8O�PObOMO�OqO�O �O�O�O�O_�OO L_#_5_�_Y_k_�_�_ �_�_ o�_�_6ooo loCoUogo�o�o�o�o �o�o �o	h�O �w�����
� �.�	__I'�1_� q��������ˏݏ� ��%�r�I�[���� ������ǟٟ&���� \�3�E�W����ȯ�� �ׯ�"��F�1�j� E�s�����m������� ѿ�0���f�=�O� a�sυϗ��ϻ���� ����'�9�Kߘ�o� ������[����(�� L�7�p��m��� ��������$����� l�C�U���y������� ���� ��	V-? �cu����
 ��@+dO�s ��������*/ //`/7/I/[/m// �/�/�/�/?�/�/? !?3?E?�?i?{?�?�? �?�?�?�?�?FO�jO UOgO�O�O�O�O�O�O __�'O9OO=_O_ �_s_�_�_�_�_�_�_ �_oPo'o9o�o]ooo �o�o�o�o�o�o: #5��O��� �� ��$��H�Fz��$DCSS_S�LAVE ;����w���`�_4D  �w���AR_MEN/U <w� >�؏@���� �2�^rǏ�\�n�\���SHOW� 2=w� � fr[q����Ə��� ��,�>�D�b�t��� ����ҟϯ��� �)�P�M�_�q����� ����˿ݿ���:� 7�I�[ς�|Ϧ��ϵ� ��������$�!�3�E� l�fߐύߟ߱����� �����/�V�P�z� w����������� ��@�:�d�a�s��� ��������\���*� H�N�K]o��� �����28� GYk}���� ��"�1/C/U/ g/y/�/��/�/�/� �//?-???Q?c?u? �/�?�?�?�/�??O O)O;OMO_O�?�O�O �O�?�O�?�O__%_ 7_I_pOm__�_�O�_ �O�_�_�_o!o3oZ_ Woio{o�_�o�_�o�o �o�oDo-Se �o��o�������.�=�O���CFoG >������q��dMC:�\��L%04d.'CSV\��pc����m���A ՃCH݀�z�v�w�#��q���:�J�8�7����JP�j�)�́�p+�n�RC_O�UT ?z����a�_C_F�SI ?�� |���� �@�;�M�_������� ��Я˯ݯ���%� 7�`�[�m�������� ǿ�����8�3�E� Wπ�{ύϟ������� �����/�X�S�e� wߠߛ߭߿������� �0�+�=�O�x�s�� ������������ '�P�K�]�o������� ����������(#5 Gpk}���� � �HCU g������� � //-/?/h/c/u/ �/�/�/�/�/�/�/? ?@?;?M?_?�?�?�? �?�?�?�?�?OO%O 7O`O[OmOO�O�O�O �O�O�O�O_8_3_E_ W_�_{_�_�_�_�_�_ �_ooo/oXoSoeo wo�o�o�o�o�o�o�o 0+=Oxs� �������� '�P�K�]�o������� ����ۏ���(�#�5� G�p�k�}�������ş ן �����H�C�U� g���������دӯ� �� ��-�?�h�c�u� ��������Ͽ���� �@�;�M�_ψσϕ� ������������%� 7�`�[�m�ߨߣߵ� ���������8�3�E� W��{��������� �����/�X�S�e� w��������������� 0+=Oxs� ����� 'PK]o��� �����(/#/5/ G/p/k/}/�/�/�/�/ �/ ?�/??H?C?U3��$DCS_C_�FSO ?�����1 P [?U?�?�? �?�?�?O
OO.OWO ROdOvO�O�O�O�O�O �O�O_/_*_<_N_w_ r_�_�_�_�_�_�_o oo&oOoJo\ono�o �o�o�o�o�o�o�o' "4Foj|�� �������G� B�T�f���������׏ ҏ�����,�>�g� b�t���������Ο�� ���?�:�L�^����������ϯʯܯg?C/_RPI~>�?� ;�d�_�
�}?.�p���X�ݿj>SL�@�� �9�b�]�oρϪϥ� �����������:�5� G�Y߂�}ߏߡ����� �������1�Z�U� g�y���������� ��	�2�-�?�Q�z�u� ������������
 )RM_q�� �����*% 7Irm��� ��/�ϛ�,�/ W/�/{/�/�/�/�/�/ �/???/?X?S?e? w?�?�?�?�?�?�?�? O0O+O=OOOxOsO�O �O�O�O�O�O___ '_P_K_]_o_�_�_�_ �_�_�_�_�_(o#o5o Gopoko}o�o�o�o�o �o �oHCU g��������� ����NOCO�DE @������PRE_?CHK B��3��A 3��< �7��������� 	 <�����?# ۏ%�7��[�m�G�Y� ������ٟ�ş�!� ���W�i�C�����y� ïկˏ������A� S�-�_���c�u���ѿ �������=��)� sυ�_ϩϻϕ����� ���'�9���E�o�I� [ߥ߷ߑ��������� #����Y�k�E��� {����������� C�U��=�����w��� ������	����?Q +u�a���� ��);_q g�Y��S��� �%/�/[/m/G/�/ �/}/�/�/�/�/?!? �/E?W?1?c?�?�� �?�?o?�?O�?�?AO SO-OwO�OcO�O�O�O �O�O_�O+_=__I_ s_M___�_�_�_�_�_ �?�_'o9oo]oooIo �o�oo�o�o�o�o #�oGY3E�� {�����o� C�U��y���e����� ������	��-�?�� K�u�O�a�������� �͟��)��1�_�q� �}�������ݯ�ɯ �%���1�[�5�G��� ��}�ǿٿ����� ��E�W�1�{ύ�G�u� ���ϯ������/�A� �-�w߉�c߭߿ߙ� ��������+�=��a� s�M���ϑ����� ���'��3�]�7�I� ������������� ����GY3}�i �������� C/y�e�� �����-/?// c/u/O/�/�/�/�/�/ �/�/?)?�?_?q? K?�?�?�?�?�?�?�? O%O�?IO[O5OO�O kO}O�O�O�O�O_�O 3_E_;?-_{_�_'_�_ �_�_�_�_�_�_/oAo oeowoQo�o�o�o�o �o�o�o+7a W_i_��C��� ��'��K�]�7�i� ��m��ɏۏ����� ��G�!�3�}���i� ��ş������1� C��g�y�S�e����� �����ѯ�-��� c�u�O�������Ͽ� ןɿ�)�ÿM�_�9� kϕ�oρ����Ϸ�� ����I�#�5�ߑ� kߵ��ߡ������� 3�E���Q�{�U�g�� ����������/�	� �e�w�Q��������� ������+Oa �I������ �K]7� �m�����/ �5/G/!/k/}/se/ �/�/_/�/�/�/?1? ??g?y?S?�?�?�? �?�?�?�?O-OOQO cO=OoO�O�/�/�O�O {O�O_�O_M___9_ �_�_o_�_�_�_�_o o�_7oIo#oUooYo ko�o�o�o�o�o�O�o 3Ei{U�� ������/�	� S�e�?�Q�������я ㏽����O�a� ������q���͟���� ���9�K�%�W��� [�m���ɯ�����ٯ �5�+�=�k�}���� ���������տ�1� �=�g�A�Sϝϯω� ���Ͽ�������Q��c����$DCS_SGN CS�����#M��25-JUN-�24 10:34� E�06��0O9:39������ X�L��ԁ����������Дќ�M��Þ��j�����{�VERSION ���V4.2.1�0�EFLOGI�C 1DS��  	D����X�k�X�z�M�PR�OG_ENB  ���b��Л�UL�SE  ����M�_ACCLIM^�������WRSTJNT��v���w�EMO����ѷ�L��INIT� EZ�O��O�PT_SL ?	�S�1�
 	Rg575�Ӆ�74���6��7��5A��1���2��l���G�h�TO  t���.H�]V?�DEX��d�����FPATH ;A��A\4����HCP_CL?NTID ?+�b� l������IAG_GRP �2JS�� �a[�D��  D�� D�  B�  B��@ff��/B!�@[��W�@��q��B�N��C�-Bz���Bp@e`���mp3m7 7�89012345�6�*�[��  �Ao�mAj�1AdA]��
AW|�AP���AJ-AC/A;�A4H|���@�  A��eA�A3!_A�@�@��B4�� ���t���
�u���ApffAj��yAeK�A_�AY��AS� �MC�AF��A@ �O�+/=/O$O�xc K�w(@�X?�8��@��y��/�/�/�/�/8�;�d�2�5?@~f�f@x1'@q���@kC�@d��D@]��@Vv��6?H?Z?l?~?8s��0l��@e�@^��@W\)�@O��@H�0?�<@7K�@.V��?�?�?�?
O8S�@M00G<@A���@<1@5���@/l�@(�w�@!�0�\NO `OrO�O�Ox'g�L_K� ;_�_�__g_�_�_�_ �_o�_�_�_YokoIo �o�o+o�oX�"� �2�17A�@J>���R
q?�33?Y���r��J7�'Ŭ2q63p4��F>r��LJ@��p�Zr�
=@�@�Q�jqZ��@G Ah�@��@��T= c<���]>*�H>�V>�3�>����J<���<��p�q�x��� ��?� �C�  �<(�U�� 4Vr�33��@
���A@��?R�oD��m R�x���Q��t����Z��Џ��؏�,��i?��7N�>�(�>��@Z�=���J�7�G�v�G�J�B��E�����a��@ǐ@����@��@Q��?L �����I�P���&���'��@�K����A�g�q�PC�  C���Cuy�
����ʯ ?յ�V�?�)�Yӌ�5��V���2����=�Y�K�)�Cz�C�8�D��p �e���P6���Z��v����*
��3��6C �F�ǿB���ֿ����E�T���� =�2�������=��^>��&$
�Iϗ�C�T_CONFIG� K3����eg��ST�BF_TTS��
@����"�������{��MAU���MS�W_CF��L � K �OCVIE�W	�MI�U�� ��߭߿��������� ���0�B�T�f�x�� ������������� ,�>�P�b�t������ ����������(: L^p���� �� �6HZ l~�����X�/��RCB�N��!�X.F/{/j/�/��/�/�/�/��SBL�_FAULT �O9*^�1GPMS�K��7��TDIAOG P��U�����qUD1�: 6789012345q2�q���%P�ϭ?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O �a6�I'��
�?_��TREC	PJ?\:
j4\_�7u[ �?�_�_�_�_�_�_o o(o:oLo^opo�o�o��o�o�O�O_ _�U�MP_OPTIO1N��>qTRB���:9;uPME��.�Y_TEMP  È�3B����p�A�pytUNI�'��ŏq6�YN_B�RK Qt�_�EDITOR q&qh��r_2PENT 1�R9)  ,&�COLOCA_�BARRA_�pN�O &p5� &�MAIN '�ES�TEIRA2���&PEG%�W����& �bpA_I�RVIS$r�� �&PICKUP*��M�P�p 
���&-BCKE�DT- ُ�S�EGU*�'��=� �&SUMIRG_SE����T��F+�DA_PRE'NSAg���Є���0� A����Ё1?_PLACE0���&
x�-�,�Ᶎ��&T�'���� v�у'�C���ޒ,����o�U���'����\�����G� ���6�<Ĉ��BASE��=���/t�����EMG?DI_STA�u~���q�uNC_INF�O 1SI��b�������Կⷮ���;1TI� ��o#���G�d�o}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������Hu� �2�D� R�j�R�x������ ��������,�>�P� b�t������������� Z��#5Ga�k }������� 1CUgy� �������	// -/?/Yc/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?��?O%O7OQ/GO mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�?Oo o/o�_[Oeowo�o�o �o�o�o�o�o+ =Oas���� ��_�_��'�9�So ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�K�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�C� 5�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������ ���!�;�M�W�i�{� ������������� �/�A�S�e�w����� ����������+ E�Oas���� ���'9K ]o����1�� ��/#/=G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?��?�?	OO 5/?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�? �_�_oo-O#oIo[o moo�o�o�o�o�o�o �o!3EWi{ ����_�_��� �7oA�S�e�w����� ����я�����+� =�O�a�s�������� �ߟ���/�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������͟׿��� �'�1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ſ���������;� M�_�q������� ������%�7�I�[� m�������߯����� ���)�3EWi{ ������� /ASew�� �������/!+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?/��?�? �?�?/#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�?�_�_�_�_Oo -o?oQocouo�o�o�o �o�o�o�o); M_q���_�� ��	o�%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ����ß՟矝�� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߩ���������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u����߫� ����������); M_q����� ��%7I[ m�������� /!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�� �?�?�?�?�OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�?�?�_�_�_�_ �?�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy�_ �����_�	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q��y�����˟ �۟��%�7�I�[� m��������ǯٯ� ���!�3�E�W�i���� �$ENETM�ODE 1U���  
��������»���RROR_PRO/G %��%������TABLE  ���Q�c�u�����SEV_NU�M ��  �������_AU�TO_ENB  q̵��ݴ_NO��� V�������  *��������������+���(�<:���FLTR���ƇHIS�Ð�����_�ALM 1W��� ����̍�+ ;���������0�?߹_����  �����²u꒰TCP_�VER !��!���@�$EXTLO�G_REQv������SIZ����SkTK�������TOL  ��D�z~��A ��_BWDU�*�Z�V�ǲv?�DID� X敇Z�����[�S�TEPl�~�����O�P_DO���FA�CTORY_TU�Nv�d��DR_G�RP 1Y��`�d� 	p�.° ��*u���R�HB ��2 ���� �e9 ����bt� A��5�BB��\B-ܵAލ�B~A���@��-A����B&�A����A��BX�� ����
C.�gR  >�Β�A�T@ICm�u��
 J)�q�����AZR����a[ /�$/�B��  F!A�  �@�33R"�33.�UUTn*@P  �/ȷ>u.�>*���<��ǊE�� F@ �"�5W�%�J���NJk�I'P�KHu��IP��sF!���?��  ?�/9�<�9�89�6C'6<,�5����Zk���̅���F��� y�U��t{G �FEAT?URE Z�V��ƱHan�dlingToo�l �5��En�glish Di�ctionary��74D St�0a�rd�6�5Anal?og I/O�7�7�gle Shif�t Outo So�ftware U�pdate%Ima�tic Back�up�9SAground Edit�0~�7Camera�0�F�?CnrRnd�ImXC�Lommo�n calib �UI�C�FnqA�@M�onitor�Kt�r�0Reliab<@�8DHCP�IZ�ata Acqu�is�CYiagn�osOA�1[ocu�ment Vie�we�BWual �Check Sa�fety�A�6ha�nced�F�:�Us�nPFr�@�7xt.� DIO �@fi�RT�Wend�PErEr�@LQR�]�Ws�Y�r�0�P E�:FCTN Menu�P�v S8gTP In�'`facNe�5Gi�gE`nrej@p Mask Exc�P�g�WHT^`Pro�xy SvoT�fi�gh-Spe�PS�ki�D�eJP�Pmm�unicN@ons�hurE`'`_�1ab�connect �2xncr``st#ru�2z>peeQP�JQU�4KAREL Cmd. L�`�ua�husRun-;Ti�PEnvkx(`�el +R@sP@S�/W�7Licen�se�Sn\�PBoo�k(System�)�:MACROs�,�b/Offse�@�uH�P8@_�pM�R�@�BP^Mech/Stop�at.p6R"�ui�RKj�x�P�0�P@)�od@wit#ch��>�EQ.����OptmЏ>��`f�iln\=�gw�uulti-T�`tC�9PCM funHw�F�o3T�R?�f�Re�gi�pr�`I�ri�gPFV����0Num� Selb����P Adju�`���J�tatu��
�iZ��5RDM Rob�ot�0scove��1F�ea7��PFreq Anly�g'Rem`��Qn�7F�>R�Servo�P��~�8SNPX b�rvNSN^`ClifQ<ɮBLibr�3鯢�0 q�����o�ptE`ssag?��4��a -C��;��/I_m>B�MILIBk�E�?P Firm6BU��PEcAcck@sKT�PTX_C�eln����F��1�V�or�qu@imulah�A�A�u��Pa�q�U�j@�Ã&�`ev�.B�.@riP޿�USB port- �@iP�PagP��?R EVNT�ϗ�nexcept�P`��t��ſX�]VC�Ar�b�bf�V2PҦ�h$����SܠSCص�V�SGEk�a�UI~�;Web Pl!� �ާ��Խ`�TeQf�ZDT Appl��d�:�ƺ� �Gri=dV�play�R�WD4�R
�.�:n�EQ�+��r-10iA/�7L*��1Grapghic���5dv�S7DCSJ�ck�q�5�larm Cau�se/��ed�8A�scii�a��LosadnP�Upl,�2�Ol�0�AGu�6N�`���yFyc@�r��0���PV��Jo��m� c�R���c���m�./�����Q�2*u:e�RAJ��P�ٶ4eqiqnL����8NRT����9On�0e He�l�HJ�`oI�alletiz?�H������_�tr�[ROS GEth�q��T@e�װ��!�n�%�2D�tP�kg&Up9g~�(2DV-�3D Tri-jQ:EAưDef.qEBa)pdei���, �bImπF�fЎ�nsp.q=�46�4MB DRAM�Z,#FRO5/@e3ll�<�Mshf!r/"�'c%3@pLƖ,ty@s˒xG��m��.[�� ��BUp���Q�B�=mai�P�߫�]Q����@q6wl!u���^`�xR�?eL� Sup������0�P�`cr��@�R����b䚮�pr1uest�rt~QQ��ߋ�L!�4O��q$�K���l Bui7�n���APLCOO�EV�l%��CGU�OCR�G�O��DR��O
TL�S_��BU/_��K��qN_d�TA�OxVB��_�W�ܑZ���_TC�B�_�V�_�W���WF +o�V�O�W._�W�ņoTEH�o�f�O�gt&�oTEj�xVF�_w�_xVGoTwBTw~o2xVH�xVIA��vL�xVLN�yUMz �bo�f_xVN�xV!P���^xVR&xV!S��܇ʏ��W���v���VGF:�L�P2_h��h�V�h��_g�D��h�FFoh���g�RD�� TUT&��01:�L�2V�L��TBGG��v�ra�in�UI��
%HsMI���pon��m�f�"�F�>&KAREL9� ��TPj��<6 SW�IMESTڢF0O�<5�
"a�X�j��� ����ͿĿֿ���'� �0�]�T�fϓϊϜ� ����������#��,� Y�P�bߏ߆ߘ��߼� ��������(�U�L� ^����������� ����$�Q�H�Z��� ~�������������  MDV�z� �����
 I@Rv��� ���///E/</ N/{/r/�/�/�/�/�/ �/???A?8?J?w? n?�?�?�?�?�?�?O �?O=O4OFOsOjO|O �O�O�O�O�O_�O_ 9_0_B_o_f_x_�_�_ �_�_�_�_�_o5o,o >okoboto�o�o�o�o �o�o�o1(:g ^p������ � �-�$�6�c�Z�l� ��������Ə���� )� �2�_�V�h����� ��������%�� .�[�R�d��������� ������!��*�W� N�`������������ ޿���&�S�J�\� �πϒϤ϶������� ��"�O�F�X߅�|� �ߠ߲��������� �K�B�T��x��� �����������G� >�P�}�t��������� ����C:L yp������ 	 ?6Hul ~�����/� /;/2/D/q/h/z/�/ �/�/�/�/?�/
?7? .?@?m?d?v?�?�?�? �?�?�?�?O3O*O<O iO`OrO�O�O�O�O�O �O�O_/_&_8_e_\_ n_�_�_�_�_�_�_�_ �_+o"o4oaoXojo|o �o�o�o�o�o�o�o' 0]Tfx�� �����#��,� Y�P�b�t��������� ������(�U�L� ^�p����������ܟ ���$�Q�H�Z�l� ~��������د���� �M�D�V�h����  H55�2}���21��R7�8��50��J61�4��ATUPͶ5�45͸6��VCA�M��CRI�UI�Fͷ28	�NREv��52��R63���SCH��DOCV�]�CSU��869zͷ0ضEIOC9��4��R69��ES�ET���J7��R{68��MASK���PRXY!�7��OCO��3帨���̸m3�J6˸53���H2�LCH��OP�LG�0�MHCuR��S{�MCS��0��55ضMDS�W���OP�MP�R�M�@�0̶PCM �R0���ض�ж@�51�51<�0n�PRS��69��FRD�FREQn��MCN��93̶�SNBAE�3�SH�LB��M��M���2�̶HTC�TMI�L����TPA��T7PTX��EL�����8������J95n,�TUT�95�wUEV��UEC��wUFR�VCC���O��VIP�CS�C,�CSG8�r�IWEB�HTTf�R6C�N�CG{IG��IPGS)�RC�DG�H7u7��6ضR85�ƷR66�R7��Rn:�R530�680�I2�q�J��H�6<�E6,�RJح�0�4��6o64\�5�N�VD��R6��R8�4Tg����8�9�0\���J93�91Đ 7+���,�D0:oF�CLI����CMS�� �ST�Y��TO�q���7v�NN�ORS�ֱJ% ��j�OL(E�ND��L��Sf(F;VR��V3D���wPBV,�APL��wAPV�CCG䶷CCR|�CD��C�DL@CSBt�C�SK��CT�CT!BL9��U0,(C��y0L8C��TC �y0�'�TC(7TC��CT1E\��07TEh��0V��TFd8F,(GL8)GI�8H�8I��E@\�87�CTM,(M�8UM@8N�8PHHPL8YRd8(TSd8W�In@VGF�GP2���P2���@�H{7VP�D�HF �VPSGVPR�&VT��YP���VTB7Vs�IHb��VI aH'VK��=VGene���� �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=?�O?a?s?�?  H55hT�1�1�[U�3R78�<50ޭ9J614�9AT�U�T�4545�<6έ9VCA�D�3CR�I,KUI8T�528n-JNRE�:52JwR63�;SCH�9/DOCV�JCU�4�869�;0�:EI�O�TsE4�:R69�JESET�;KJ�7KR68�JMA{SK�9PRXYML]7�:OCO\3�<h�J)P�<3|ZJ6�<�53�JH�\LCH^\ZOPLG�;0�Z�MHCR]ZSkMkCS�<0,[55�:�MDSW}k�[OP��[MPR�Z�@�\0n�:PCMLJR0�k�)P�:)`�[51K5u1|0JPRS[�69|ZFRD<JFwREQ�:MCN�:{93�:SNBA}K^�[SHLB�zM�{t�@ll2�:HTC�:�TMIL�<�JTP�A�JTPTX�EL�z)`�K8�;�0�JwJ95\JTUT�[�95|ZUEVZU�EC\ZUFR<JV�CC��O<jVIP�,�CSC\�CSGtlJ�@I�9WEB�:7HTT�:R6{L���CG{�IG[�IP�GS��RC,�DG��[H77�<6�:R�85�JR66JRu7[R|R53{K68|2�Z�@Jml*,|6|6\JR�\	Pj|4L�6�64���5�kNVDZR6+kR84<���IP,��8��90���KJ9&�\91��̫7[KIP�\JD0�F��CL9I�lKCMS�J9�n�:STY,�TO�:��@�K7�LNN|ZO�RS<jJ��MZZ|O]LK�END�:L��S��FVR�JV3�D,�KKPBV\�A�PL�JAPV�ZC�CG�:CCRjC�D�CDL̚CS�B�JCSK�jCTK�CTB��\���\��C�z���CL�TC�LJ�l�TC��TC�ZCTE�J��|�T�E�J��<�TF��FJ\�G��G��l�Hl��I�z)�l�k�CTM�\�M\�M��Nl�P�,�P��R��;�TSr��W��̚VGF��P2��P2�z ��VPDFLJV�P;�VPR��VT��;� �JVTB��V�KIH�VِM�<��VK,�V{�Gene�8�83EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{?��7�0STD~�4LANG�4 �9�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� ��2�D�V�RBT�6OPTNm�������� Ǐُ����!�3�E� W�i�{�������ß�5DPN�4����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}�x�ߡ߳�ted �4 �8��������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������@��ǯٯ�������*�<�N�`�r���9�9���$FEAT�_ADD ?	��������  	��ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu�����DEMO Z��?   ���} ��'��0�]�T�f� �������������� #��,�Y�P�b����� ������������ (�U�L�^��������� ���ܯ���$�Q� H�Z���~�������� ؿ��� �M�D�V� ��zόϦϰ������� �
��I�@�R��v� �ߢ߬��������� �E�<�N�{�r��� �����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo~o �o�o�o�o�o�o�o! *WN`z�� �������&� S�J�\�v��������� �ڏ���"�O�F� X�r�|�������ߟ֟ ����K�B�T�n� x�������ۯү�� ��G�>�P�j�t��� ����׿ο���� C�:�L�f�pϝϔϦ� ������	� ��?�6� H�b�lߙߐߢ����� ������;�2�D�^� h����������� ��
�7�.�@�Z�d��� �������������� 3*<V`��� �����/& 8R\����� ����+/"/4/N/ X/�/|/�/�/�/�/�/ �/�/'??0?J?T?�? x?�?�?�?�?�?�?�? #OO,OFOPO}OtO�O �O�O�O�O�O�O__ (_B_L_y_p_�_�_�_ �_�_�_�_oo$o>o Houolo~o�o�o�o�o �o�o :Dq hz������ �
��6�@�m�d�v� ������ُЏ��� �2�<�i�`�r����� ��՟̟ޟ���.� 8�e�\�n�������ѯ ȯگ����*�4�a� X�j�������ͿĿֿ ����&�0�]�T�f� �ϊϜ����������� �"�,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/
??A? 8?J?w?n?�?�?�?�? �?�?�?OO=O4OFO sOjO|O�O�O�O�O�O �O__9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿����&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t����������   ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�����y  �x�q��� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p��P����q�p�x ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p���������������$F�EAT_DEMO�IN  ��� �����IND�EX���I�LECOMP �[���B���8 SETU�P2 \B~L�  N w�5_AP2BCK� 1]B	  #�)����%����E �	���5 �Y�f��B ��x/�1/C/� g/��/�/,/�/P/�/ t/�/?�/??�/c?u? ?�?(?�?�?^?�?�? O)O�?MO�?qO O~O �O6O�OZO�O_�O%_ �OI_[_�O__�_�_ D_�_h_�_�_
o3o�_ Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0����ׯQ	� P� 2>� *.VRޯ(���*+�Q���W�{��e��PC������OFR6:��ؾg�����T   �2�����\� ��d�*.F��ϕ�	ó����qo�ߓ�STM� 9���ư%�d��ψ���HU߻�Jש�f�x���GIF�A�L��-����ߑ��JPG ����Lձ�n�����#JS�H�����6����%
JavaS�criptt���C�Se���Kֹ�v� %�Cascadi�ng Style Sheets���j�
ARGNAMOE.DT'��OЁ\;��[�k|(>k DISP*rU�Oп��� �
�TPEINS.X3ML/�:\C�cCustom Toolbar���	PASSWOR�D���FRS:�\�� %Pa�ssword Config/c�Q/ �J/�/���/:/�/�/ p/?�/)?;?�/_?�/ �??$?�?H?�?l?�? O�?7O�?[OmO�?�O  O�O�OVO�OzO_�O �OE_�Oi_�Ob_�_._ �_R_�_�_�_o�_Ao So�_woo�o*o<o�o `o�o�o�o+�oO�o s��8��n ��'���]���� �z���F�ۏj���� ��5�ďY�k������ ��B�T��x����� C�ҟg�������,��� P���������?�ί �u����(���Ͽ^� 󿂿�)ϸ�M�ܿq� ��ϧ�6���Z�l�� ��%ߴ��[����� �ߵ�D���h����� 3���W����ߍ��� @����v����/�A� ��e������*���N� ��r�����=��6 s�&��\� �'�K�o� �4�X��� #/�G/Y/�}//�/ �/B/�/f/�/�/�/1? �/U?�/N?�??�?>? �?�?t?	O�?-O?O�?�cO�?�OO(O�O�F��$FILE_DG�BCK 1]����@��� < �)
S�UMMARY.DyG�OsLMD:�O�;_@Diag� Summary�<_IJ
CONSLOG1__&Q_�_NQ�Console� log�_HK	T�PACCN�_o%�o?oJUTP A�ccountin��_IJFR6:I�PKDMP.ZI	PsowH
�o�oKU[`�Exceptio�n�oyk'PMEMCHECK5o�_*_K��QMemory� DataL�F�4l�)6qRIP�E�_$6�Zs%��q Packe�t L�_�DL�$y�	r�qSTAT����S� %~�rStatusT��	FTP���:����Vw�Qmmen�t TBD؏� �>I)ETHERNE���
q�[��NQEthern��p�Pfigura��oODDCSVRAF̏��ďݟd���� verify �all��{D�.���DIFF՟��͟xb��s��diffd���
q��CHG01 Y�@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ��VTRNDIAG.LS�̿޿s�^q=3� Ope���q� SQnostic��w��)VD;EV7�DATt�Q�xc�u�g�Vis��?Device�Ϫ�IMG7ºo����y�z�s�Imag�n��UP��ES��~T�FRS:\��� �OQUpdates List ��IJg�FLEXEVENQ�X�j߃�f��F� UIF E�v���B,�s��)
PSRBWLOD.CM��sL�������PPS_RO�BOWEL��GL�o�GRAPHIC�S4Dy�b�t���%4D Gra�phics Fi�leu��AOɿ��rGIG���u�
>YvGigE�ة�~�BN�? )��HADOW������\sShadow Chang���vbQRCMERR�n�\s�� CFG Er�ror�tail�� MA��C?MSGLIB� �"^o� ���T�)�ZD�����/XwZD�6 ad�HPNOTI���
/�/Zu�Notific8��H/��AGUO�/ yO?�O'?P?OOt?? �?�?9?�?]?�?O�? (O�?LO^O�?�OO�O 5O�O�OkO _�O$_6_ �OZ_�O~_�__�_C_ �_�_y_o�_2o�_?o ho�_�oo�o�oQo�o uo
�o@�odv �)�M��� ��<�N��r���� ��7�̏[������&� ��J�ُW������3� ȟڟi�����"�4�ß X��|������A�֯ e�����0���T�f� ���������O��s� �ϩ�>�Ϳb��o� ��'ϼ�K����ρ�� ��:�L���p��ϔߦ� 5���Y���}���$�� H���l�~���1��� ��g���� �2���V� ��z�	�����?���c� ��
��.��Rd�� ���M�q �<�`��� %�I��/� 8/J/�n/��/!/�/ �/W/�/{/?"?�/F? �/j?|??�?/?�?�?��$FILE_F�RSPRT  ����0�����8MDON�LY 1]�5�0� 
 �)M�D:_VDAEX?TP.ZZZ�?�?�_OnK6%N�O Back f�ile 9O�4S�6Pe?�OOO�O�?�O __?>_�Ob_t__�_ '_�_�_]_�_�_o(o �_Lo�_po�_}o�o5o �oYo�o �o$�oH Z�o~��C� g��	�2��V�� z������?�ԏ�u��
���.�@��4VIS�BCKHA&C*�.VDA�����F�R:\Z�ION\�DATA\v�����Vision VD�B��ŏ��� '�5��Y��j���� ��B�ׯ�x����1� ��үg�������X��� P��t���Ϫ�?�ο c�u�ϙ�(Ͻ�L�^� �ς��)���M���q�  ߂ߧ�6���Z���� ��%��I�������:�LUI_CONF�IG ^�5|m��� $ h�F{�5������)�;�I���|xq�s��� ��������a���  $6��Gl~�� �K��� 2 �Vhz���G ���
//./�R/ d/v/�/�/�/C/�/�/ �/??*?�/N?`?r? �?�?�???�?�?�?O O&O�?JO\OnO�O�O )O�O�O�O�O�O_�O 4_F_X_j_|_�_%_�_ �_�_�_�_o�_0oBo Tofoxo�o!o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� �����ʏ܏��� $�6�H�Z�l������ ��Ɵ؟ꟁ�� �2� D�V�h���������¯ ԯ�}�
��.�@�R� d�����������п� y���*�<�N�`��� �ϖϨϺ�����u�� �&�8�J���[߀ߒ� �߶���_������"� 4�F���j�|���� ��[�������0�B� ��f�x���������W� ����,>��b t����O���(:�  �xFS�$FL�UI_DATA �_������uRESULT 2`��� �T��/wizard�/guided/�steps/Expertb��/ /+/=/O/a/s/�/�/��*�Conti�nue with{ G�ance�/ �/�/??(?:?L?^?�p?�?�?�? T-�U��90 �`� �?���9��ps�?0OBOTOfOxO �O�O�O�O�O�O�O�  �_/_A_S_e_w_�_ �_�_�_�_�_�_n�?��?�?�<Frip �Oo�o�o�o�o�o �o�o!3E_i {������� ��/�A�S�o$on��HoAO�TimeUS/DST[� �����+�=�O�a��s������'Enabl�/˟ݟ��� %�7�I�[�m������T�?{�ݯ����Æ24Ώ3�E�W�i� {�������ÿտ翦� ���/�A�S�e�wω� �ϭϿ������ϴ�Ư�د� G��Region�χߙ߽߫� ��������)�;�+�America sou�������������)�;��?�y��#߅�G�Y��ditorL������� #5GYk}��+� Touch P�anel �� (�recommen�)���*�<N`r��U���e�w��������accesd�./@/R/d/ v/�/�/�/�/�/�/Q|�Connect� to Network�/(?:?L?^? p?�?�?�?�?�?�?�?
Y���������!/��Introducts߆O�O�O �O�O�O�O__(_:_ U^_p_�_�_�_�_�_��_�_ oo$o6oHo e�Oeo?O�X_�o �o�o�o'9K ]o��R_��� ���#�5�G�Y�k��}�����h`�ooj }oߏ�o��*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ쯫� ��Ϗ1��X�j�|��� ����Ŀֿ����� 0��A�f�xϊϜϮ� ����������,�>� ��_�!���E��߼��� ������(�:�L�^� p���߸�������  ��$�6�H�Z�l�~� ��O߱�s�������  2DVhz�� ������
. @Rdv���� ����/��'/��� `/r/�/�/�/�/�/�/ �/??&?8?�\?n? �?�?�?�?�?�?�?�? O"O4O�UO/yO�O O?�O�O�O�O�O__ 0_B_T_f_x_�_I?�_ �_�_�_�_oo,o>o Poboto�oEO�OiO�o �o�O(:L^ p�������_  ��$�6�H�Z�l�~� ������Ə؏�o�o�o �/��oV�h�z����� ��ԟ���
��.� �R�d�v��������� Я�����*���� ����C�����̿޿ ���&�8�J�\�n� ��?��϶��������� �"�4�F�X�j�|ߎ� M�_�q��ߕ����� 0�B�T�f�x���� ���������,�>� P�b�t����������� ���߱���%��L^ p�������  $��5Zl~ �������/  /2/��S/w/9�/ �/�/�/�/�/
??.? @?R?d?v?�?�/�?�? �?�?�?OO*O<ONO `OrO�OC/�Og/�O�/ �O__&_8_J_\_n_ �_�_�_�_�_�_�?�_ o"o4oFoXojo|o�o �o�o�o�o�O�o�O �O�oTfx��� ������,��_ P�b�t���������Ώ �����(��oI� m��C�����ʟܟ�  ��$�6�H�Z�l�~� =�����Ưد����  �2�D�V�h�z�9��� ]���ѿ����
��.� @�R�d�vψϚϬϾ� �Ϗ�����*�<�N� `�r߄ߖߨߺ��ߋ� տ����#��J�\�n� ������������� �"���F�X�j�|��� ������������ ������u7�� ����,> Pbt3����� ��//(/:/L/^/ p/�/ASe�/��/  ??$?6?H?Z?l?~? �?�?�?�?��?�?O  O2ODOVOhOzO�O�O �O�O�O�/�/�/_�/ @_R_d_v_�_�_�_�_ �_�_�_oo�?)oNo `oro�o�o�o�o�o�o �o&�OG	_k -_������� �"�4�F�X�j�|�� ����ď֏����� 0�B�T�f�x�7��[ �������,�>� P�b�t���������ί �����(�:�L�^� p���������ʿ��� ���џӿH�Z�l�~� �Ϣϴ����������  �߯D�V�h�zߌߞ� ����������
��ۿ =���a�s�7ߚ��� ��������*�<�N� `�r�1ߖ��������� ��&8J\n -�w�Q������ "4FXj|� �������// 0/B/T/f/x/�/�/�/ �/���/?�>? P?b?t?�?�?�?�?�? �?�?OO�:OLO^O pO�O�O�O�O�O�O�O  __�/�/�/?i_+? �_�_�_�_�_�_�_o  o2oDoVoho'O�o�o �o�o�o�o�o
. @Rdv5_G_Y_� }_����*�<�N� `�r���������yoޏ ����&�8�J�\�n� ��������ȟ��� ��4�F�X�j�|��� ����į֯����ˏ �B�T�f�x������� ��ҿ�����ٟ;� ��_�!��ϘϪϼ��� ������(�:�L�^� p߁ϔߦ߸�������  ��$�6�H�Z�l�+� ��Oϱ�s��������  �2�D�V�h�z����� ����������
. @Rdv���� }�������<N `r������ �//��8/J/\/n/ �/�/�/�/�/�/�/�/ ?�1?�U?g?+/�? �?�?�?�?�?�?OO 0OBOTOfO%/�O�O�O �O�O�O�O__,_>_ P_b_!?k?E?�_�_{? �_�_oo(o:oLo^o po�o�o�o�owO�o�o  $6HZl~ ���s_�_�_�� �_2�D�V�h�z����� ��ԏ���
��o.� @�R�d�v��������� П�������� ]����������̯ޯ ���&�8�J�\�� ��������ȿڿ��� �"�4�F�X�j�)�;� M���q��������� 0�B�T�f�xߊߜ߮� m���������,�>� P�b�t�����{� �ϟ����(�:�L�^� p���������������  ��6HZl~ ������� ��/��S�z�� �����
//./ @/R/d/u�/�/�/�/ �/�/�/??*?<?N? `?�?C�?g�?�? �?OO&O8OJO\OnO �O�O�O�Ou/�O�O�O _"_4_F_X_j_|_�_ �_�_q?�_�?�_�?�_ 0oBoTofoxo�o�o�o �o�o�o�o�O,> Pbt����� ����_%��_I�[� ��������ʏ܏�  ��$�6�H�Z�~� ������Ɵ؟����  �2�D�V��_�9��� ��o�ԯ���
��.� @�R�d�v�������k� п�����*�<�N� `�rτϖϨ�g����� ������&�8�J�\�n� �ߒߤ߶��������� ��"�4�F�X�j�|�� �������������� ����Q��x������� ��������,> P�t����� ��(:L^ �/�A��e����  //$/6/H/Z/l/~/ �/�/a�/�/�/�/?  ?2?D?V?h?z?�?�? �?o���?�O.O @OROdOvO�O�O�O�O �O�O�O�/_*_<_N_ `_r_�_�_�_�_�_�_ �_o�?#o�?Go	Ono �o�o�o�o�o�o�o�o "4FXio|� �������� 0�B�T�ou�7o��[o ��ҏ�����,�>� P�b�t�������iΟ �����(�:�L�^� p�������e�ǯ��� ����$�6�H�Z�l�~� ������ƿؿ�����  �2�D�V�h�zόϞ� ���������Ϸ��ۯ =�O��v߈ߚ߬߾� ��������*�<�N� �r��������� ����&�8�J�	�S� -�w���c��������� "4FXj|� �_����� 0BTfx��[� �������/,/>/ P/b/t/�/�/�/�/�/ �/�/�?(?:?L?^? p?�?�?�?�?�?�?�? ����EO/lO~O �O�O�O�O�O�O�O_  _2_D_?h_z_�_�_ �_�_�_�_�_
oo.o @oRoO#O5O�oYO�o �o�o�o*<N `r��U_��� ���&�8�J�\�n� ������couo�o鏫o �"�4�F�X�j�|��� ����ğ֟蟧��� 0�B�T�f�x������� ��ү������ُ;� ��b�t���������ο ����(�:�L�]� pςϔϦϸ�������  ��$�6�H��i�+� ��O������������  �2�D�V�h�z��� ]���������
��.� @�R�d�v�����Y߻� }����ߣ�*<N `r������ ���&8J\n ��������� /��1/C/j/|/�/ �/�/�/�/�/�/?? 0?B?f?x?�?�?�? �?�?�?�?OO,O>O �G/!/kO�OW/�O�O �O�O__(_:_L_^_ p_�_�_S?�_�_�_�_  oo$o6oHoZolo~o �oOO�OsO�o�o�O  2DVhz�� �����_
��.� @�R�d�v��������� Џ⏡o�o�o�o9��o `�r���������̟ޟ ���&�8��\�n� ��������ȯگ��� �"�4�F���)��� M���Ŀֿ����� 0�B�T�f�xϊ�I��� ����������,�>� P�b�t߆ߘ�W�i�{� �ߟ���(�:�L�^� p���������� ���$�6�H�Z�l�~� �������������� ��/��Vhz�� �����
. @Qdv���� ���//*/</�� ]/�/C�/�/�/�/ �/??&?8?J?\?n? �?�?Q�?�?�?�?�? O"O4OFOXOjO|O�O M/�Oq/�O�/�O__ 0_B_T_f_x_�_�_�_ �_�_�_�?oo,o>o Poboto�o�o�o�o�o �o�O�O%7�_^ p�������  ��$�6��_Z�l�~� ������Ə؏����  �2��o;_���K ��ԟ���
��.� @�R�d�v���G����� Я�����*�<�N� `�r���C���g���ۿ ����&�8�J�\�n� �ϒϤ϶����ϙ��� �"�4�F�X�j�|ߎ� �߲����ߕ�����˿ -��T�f�x���� ����������,��� P�b�t����������� ����(:��� �A�����  $6HZl~ =�������/  /2/D/V/h/z/�/K ]o�/��/
??.? @?R?d?v?�?�?�?�? �?��?OO*O<ONO `OrO�O�O�O�O�O�O �/�O�/#_�/J_\_n_ �_�_�_�_�_�_�_�_ o"o4oE_Xojo|o�o �o�o�o�o�o�o 0�OQ_u7_�� ������,�>� P�b�t���Eo����Ώ �����(�:�L�^� p���A��eǟ���  ��$�6�H�Z�l�~� ������Ưد�����  �2�D�V�h�z����� ��¿Կ�������+� �R�d�vψϚϬϾ� ��������*��N� `�r߄ߖߨߺ����� ����&��/�	�S� }�?Ϥ���������� �"�4�F�X�j�|�;� ������������ 0BTfx7��[� �����,> Pbt����� ���//(/:/L/^/ p/�/�/�/�/�/�� ��!?�H?Z?l?~? �?�?�?�?�?�?�?O  O�DOVOhOzO�O�O �O�O�O�O�O
__._ �/�/?s_5?�_�_�_ �_�_�_oo*o<oNo `oro1O�o�o�o�o�o �o&8J\n �?_Q_c_��_�� �"�4�F�X�j�|��� ����ď�oՏ���� 0�B�T�f�x������� ��ҟ����>� P�b�t���������ί ����(�9�L�^� p���������ʿܿ�  ��$��E��i�+� �Ϣϴ����������  �2�D�V�h�z�9��� ����������
��.� @�R�d�v�5ϗ�Yϻ� }������*�<�N� `�r������������� ��&8J\n ���������� ��FXj|� ������// ��B/T/f/x/�/�/�/ �/�/�/�/??�# �G?q?3�?�?�?�? �?�?OO(O:OLO^O pO//�O�O�O�O�O�O  __$_6_H_Z_l_+? u?O?�_�_�?�_�_o  o2oDoVohozo�o�o �o�o�O�o�o
. @Rdv���� }_�_�_�_��_<�N� `�r���������̏ޏ �����o8�J�\�n� ��������ȟڟ��� �"����g�)��� ����į֯����� 0�B�T�f�%������� ��ҿ�����,�>� P�b�t�3�E�W���{� ������(�:�L�^� p߂ߔߦ߸�w�����  ��$�6�H�Z�l�~� ����������� ��2�D�V�h�z����� ����������
-� @Rdv���� �����9�� ]������� �//&/8/J/\/n/ -�/�/�/�/�/�/�/ ?"?4?F?X?j?)�? M�?qs?�?�?OO 0OBOTOfOxO�O�O�O �O/�O�O__,_>_ P_b_t_�_�_�_�_{? �_�?oo�O:oLo^o po�o�o�o�o�o�o�o  �O6HZl~ �������� �_o�_;�e�'o���� ��ԏ���
��.� @�R�d�#�������� П�����*�<�N� `��i�C�����y�ޯ ���&�8�J�\�n� ��������u�ڿ��� �"�4�F�X�j�|ώ� �ϲ�q�������	�˯ 0�B�T�f�xߊߜ߮� ���������ǿ,�>� P�b�t������� ������������[� ߂�������������  $6HZ�~ �������  2DVh'�9�K� �o����
//./ @/R/d/v/�/�/�/k �/�/�/??*?<?N? `?r?�?�?�?�?y�? ��?�&O8OJO\OnO �O�O�O�O�O�O�O�O _!O4_F_X_j_|_�_ �_�_�_�_�_�_o�? -o�?QoOxo�o�o�o �o�o�o�o,> Pb!_����� ����(�:�L�^� o�Ao��eog�܏�  ��$�6�H�Z�l�~� ������s؟����  �2�D�V�h�z����� ��o�ѯ�����˟.� @�R�d�v��������� п����ş*�<�N� `�rτϖϨϺ����� �������/�Y�� �ߒߤ߶��������� �"�4�F�X��|�� ������������� 0�B�T��]�7߁��� m�������,> Pbt���i�� ��(:L^ p���e�w����� ���$/6/H/Z/l/~/ �/�/�/�/�/�/�/�  ?2?D?V?h?z?�?�? �?�?�?�?�?
O�� �OO/vO�O�O�O�O �O�O�O__*_<_N_ ?r_�_�_�_�_�_�_ �_oo&o8oJo\oO -O?O�ocO�o�o�o�o "4FXj|� �__������ 0�B�T�f�x������� moϏ�o�o�,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ���!��E��l�~� ������ƿؿ����  �2�D�V��zόϞ� ����������
��.� @�R��s�5���Y�[� ��������*�<�N� `�r����g����� ����&�8�J�\�n� ������c��������� ��"4FXj|� �������� 0BTfx��� ����������#/ M/t/�/�/�/�/�/ �/�/??(?:?L? p?�?�?�?�?�?�?�?  OO$O6OHO/Q/+/ uO�Oa/�O�O�O�O_  _2_D_V_h_z_�_�_ ]?�_�_�_�_
oo.o @oRodovo�o�oYOkO }O�O�o�O*<N `r������ ��_�&�8�J�\�n� ��������ȏڏ��� �o�o�oC�j�|��� ����ğ֟����� 0�B��f�x������� ��ү�����,�>��P��!�3������$�FMR2_GRP� 1a���� �C4 w B�[�	 [��߿�ܰE�� �F@ 5W��S�ܰJ��NJ�k�I'PKH�u��IP�sF�!���?�  �W�S�ܰ9�<9��896�C'6<,5����A�  l�Ϲ�BHٳB�հ�����@�33�33S�۴��ܰ/@UUT'�@��8���W�>u.�>*���<����=�[�B=���=�|	<�K�<�q�=�mo����8�x	7�H<8�^6�Hc7��x?� ���������"��F��X���_CFG =b»T Q������X�NO ^º
F0�� ���W�RM_CHKTYP  ��[�ʰ�̰����ROM�_�MIN�[����9����X��SSB�h�c�� ݶf�[�]�����^�TP_DEF_�O�[�ʳ��I�RCOM���$�GENOVRD_�DO.�d���TH�R.� dd��_�ENB�� ��RWAVC��dO�Z�� ���Fs  �G!� GɃ��I�C�I(i J���+���%�q���� �Q�OU��j¼��8����<6�i��C�;]�[�C�  D�+��3@���B���p�.��R SMT���k_	ΰ\��$HoOSTCh�1l¹�[��d�۰ M5C[���/Z�  27.0� =1�/  e�/? ?'?9?G:�/j?|?�?�?�,Z?T3	anonymouy �?�?�	OO-O?N�/ڰRH RK�/�?�O�/�O�O�O �O_V?3_E_W_i_�O &_�?�_�_�_�_�_@O �_dOvOSo�_�Ojo�o �o�o�o_�o+ =`o�_�_���� �o&o8oJoL9��o ]�o��������oɏۏ ����4�j+�Y�k� }��������� � �T�1�C�U�g����� ������ӯ��x�>�� -�?�Q�c�����Ο�� �Ͽ����)�;� ��_�qσϕϧ�ʿ � �����%�7�~��� ��߶ϣ�������� ���Ϻ�3�E�W�i�� ���ϱ���������@� R�d�v�x�J��߉��� ���������+ =`���������:$h!ENT 1=m P!V  7 ?. c&�J�n�� �/�)/�M//q/ 4/�/X/j/�/�/�/�/ ?�/7?�/?m?0?�? T?�?x?�?�?�?O�? 3O�?WOO{O>O�ObO �O�O�O�O�O_�OA_ _e_(_:_�_^_�_�_��_�ZQUICCA0�_�_�_?od1@oo.o�od2�olo~o��o!ROUTE�R�o�o�o/!P�CJOG0!�192.168�.0.10	o�SC�AMPRT�\!�pu1yp��vRT��o��� !S�oftware �Operator? Panel�m�n��NAME �!�
!ROBO��v�S_CFG �1l�	 ��Auto-s�tarted'�FTP2��I�K 2��V�h�z������� ԟ����	���@� R�d�v���	����� ��:���)�;�M�_� &���������˿�p� ��%�7�I�[��"� 4�F�ڿ�������� !�3���W�i�{ߍߟ� ��D���������/� vψϚ�w�ߛ��Ͽ� ��������+�=�O� a�������������� ��8�J�\�n�p�]�� ��������� #5X�k}� ���0/D 1/xU/g/y/�/RH/ �/�/�/�//?�/?? Q?c?u?�?���/ ?�?:/O)O;OMO_O &?�O�O�O�O�O�?pO __%_7_I_[_�?�? �?t_�O�_O�_�_o !o3o�OWoio{o�o�_ �oDo�o�o�o�����_ERR n���-=vPDUSI�Z  �`^�P��Tt>muWRD �?΅�Q�  �guest �f������~��SCDMNGRPw 2o΅Wp���Q�`���fK�L� 	P01.�05 8�Q  � �|��  �;|��  ~z[ ���w����*���Ť�x����[ݏȏ���בPԠ�������)����D�r���؊p"*�Pl�P���Dx���dx�*�����%�_GWROU7�pLyN���	/�o���QU%P��UTu� ��TYàL}?pT�TP_AUTH �1qL{ <!iPendan���o֢!KAREL:*�������KC��ɯۯ���VISION SET�9����P�>� h��f�����������ҿ����X�CTRL rL}O�u���a
��eFF�F9E3-ϝTF�RS:DEFAU�LT��FAN�UC Web Server�ʅ�t� X���t@���1�C��U�g�;tWR_CONFIG s;�� ��=qIDL_CPU_PC����aBȠP�� BH��MIN�܅q��?GNR_IOFq{r��`Rx��NPT_S_IM_DO���STAL_SCR�N� �.�INT�PMODNTOL8Q����RTY0���8�-�\�ENBQ�-����OLNK 1tL{�p�������)�;�M���MAST�E�%���SLAV�E uL|�RA?MCACHEk�c�}O^�O_CFG�������UOC�����CMT_OP���Pz�YCL������_?ASG 1v;��q
 O�r��� ����&8pJ\W�ENUMzs5Py
��IP����RTRY_CN���M�=�zs���Tu ������w���p/��p��P_MEMB?ERS 2x;�l�k $��X"��?��Q'W/i)��RCA_�ACC 2y��  X�j� ��O��b6\�"  %��Q�&�#�#�/�!���,�$BUF0�01 2z�= �hTu0  uW0hf:4v:4�:4U�:4�:4�:4�:4��:4�:3i=0�2*�4"�42�4D�494UiA4iI4iQ4iY4Uia4ii4iq4iy4�i�4j�4j�4j#*�43�4E�4U�4A4�jI4jQ4jY4j���4��4�'�  �'�f94fejDu�jD�jD�jDQDf��jD�jD�jD�:3g��D�DDgDgZ!Dg)Dgg�Dw:4� +� �@h�4hJ�4h�4h�492$? 63:1@1ERI0ERQ0ER Y0ERa0ERi0ERq0ER y0ER�0:1�1�R�0�R �0�R�0�R�0�RBT�1 �RRT�1�RbT�1�RrT �1�R�T�1:1 Ab�T Ab@b!@b)@b JT8AbZTHAbQ@b Y@ba@bAhA:1pAub y@ub�@ub�@ubZd�A ub�@ub�@ub�@:1�A �b�@�bd�A�b*d�A �b�@�b�@ER�@�A Q@ER�TQER�T93-_ 65GSNrI2WSNrY2gS Nri2wSNry2�S���3 �S�r�2�S�r�2�S�r St�3�S�rkt�3�S�r �t�3�S�� Cc�B c�!B/c�St8CGc �ktPC_c�aBocv� qBcv��B�cv�c��C �cv��B�c���C�cƂ #��C�cƂ;��C�cNr �BsNr�tSs�Ԝ!��2{�4r�}ŋ���<����o�o��2�HIS!2}�� ܷ! 202?4-06-2���a��П���  �� 7 X��;  `�h�� ��0�B�T�f���X�cN��1O�������ɯ> � 9 �o��cP�-��$�6�H�n��mv��06���~���������Z��M 9 !�Բmv��;M �����r� +�!u�b�tφϘϪ� ���������;�M�:� L�^�p߂ߔߦ߸��� ���%��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��o��,P����o���P�����c�:�	b��d!�A� A gy�y��������	�96 a >��Q6HZlZ��l������&0@(�AѰ;: cF; �o�c�/1/C/�� ��P/�/�/�/�/�/�/ �/	??R/d/v/c?u? �?�?�?�?�?�?�?O <?N?;OMO_OqO�O�O �O�O�O�OO&O_%_ 7_I_[_m__�_�_�_ ��5p�����o$o6o����Td�Vb!� f�mczo�o�o�o�� �o�o
. �B��B��a��BrN`r �r��o������Xc�rѰk� ��� �@�R�d��O�O��� ��Џ����*�<� N�������������̟ ޟ���&�]�o�\� n���������ȯگ� ��5�G�4�F�X�j�|��������Ŀֿ�^I_�CFG 2~�[� H
Cycl�e Time��Busy�Idyl��min�=S�Up���Read(��DowG�C�X���Count�	ONum ������̸p����PROmG���U�P��)/softp�art/genl�ink?curr�ent=menu�page,1133,1�C�U�g�y��Tä�SDT_IS�OLC  �Y�� ���J23_�DSP_ENB � ��T���INC� ��ݸs��A �  ?�  =�?��<#�
���:�o �2�Dﰸq/�l���OB��C���O��ֆ�G_GROUP 1���{	!d<*�P����t�?�����pQ'�L�^�p�/� ���������\�~��G_IN_AUT�O����POSRE����KANJI_�MASK0��DR�ELMON ��[�ϸry���������f�Ã����Ӹt-��KCwL_L NUM���G$KEYLOGOGINGD�P�������LANGUA_GE �U���DEFAUgLT ��QLG������S��qx��$�8T�H  ���p'0���p;�p&�K͸u;��
�*!(UT1:\ J/ L/Y/k/}/ �/�/�/�/�/�/�/$>�(�H?�VLN_D?ISP ���P��&�$�^4OCTOL�TdDz����
�1GBOOK ��Ad4V�11�0� %O!O3OEOWOiKyM0�TËIgF	�5)�����O}���2_B�UFF 2��� ��p2O�_�2 ��6_M�R_d_�_�_�_ �_�_�_�_�_o3o*o <oNo`o�o�o�o�o��~�ADCS ��� ���L�O��+=�Oa�dIO 2���k +����������� �*�:�L�^�r����� ����ʏ܏���$��6�J�uuER_ITM��d������ǟٟ ����!�3�E�W�i� {�������ïկ���8��7x�SEVD��]t�TYP�����s������)RST�e�eSCRN_F�L 2��}��� ��/�A�S�e�w�F��TP{��b��=NGNAM��E�n�dUPSf0GI���2����_LO{AD��G %���%PICKUP�_COM��EPT�OR�ϖ�MAXU�ALRMb2�@����
K���_PRD��2  �3�AK�Ci0��qO=_'X�Ӭ��P 2��; �j*V	����
* ���4��*��'�`� 	xN��z������ �����1�C�&�g�R� ��n�����������	 ��?*cFX� ������ ;0q\��� ����/�/I/ 4/m/X/�/�/�/�/�/ �/�/�/!??E?0?i? {?^?�?�?�?�?�?�? �?OOAOSO6OwObO��OD�DBGDEF ��գѢѤO�@�_LDXDISA�����ssMEMO_{AP��E ?��
 �A�H$_6_�H_Z_l_~_�_�_K�F�RQ_CFG �����CA �G@i��S�@<��d%�\�o�_�P�Ґ�����*Z`/\b **:eb�DXo jho�F�o�o�o�o�o �o;�O��dZ�`U�y|��z,(9 �Mt���1��B� g�N���r���������̏	���?�A�IS�C 1���K` � �O�����O���O֟�����K�]�_MSTR� �3��SCD 1�]��l�� ��{�����دïկ� ��2��V�A�z�e��� ����Կ������� @�+�=�v�aϚυϾ� ����������<�'� `�K߄�oߨߓߥ��� �����&��J�5�Z� ��k���������� ����F�1�j�U��� y��������������0T?x�MK��Q�,��Q�$M�LTARM�R�:?g� ~s�@����@METPU��@l��4�ND�SP_ADCOLx�@!CMNT7 *FNSW(FSTLIxi%� �,����Q�|�*POSCF�=bPRPMV��ST51�,� 4�R#�
g!|qg% w/�'c/�/�/�/�/�/ �/?�/?G?)?;?}? _?q?�?�?�?�?�1*�SING_CHK�  {$MODA�S�e���#E�DEV 	�J	�MC:WLHSI�ZE�Ml �#ETA�SK %�J%$�12345678�9 �O�E!GTRI�G 1�,� l �Eo#_�y_S_�}�F�YP�A�u9D"CE�M_INF 1��?k`)AT?&FV0E0X_�]�)�QE0V1&�A3&B1&D2�&S0&C1S0}=�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_�_o �3o��o���o� �"�4��X��� ASe֏���C� 0���f�!���q��� ��s�䟗�����͏>� �b���s���K���w� ��ٯ�ɟ۟L��� �#�����Y�ʿ�� ����$�߿H�/�l�~� 1���U�g�y����ϯ�  �2�i�V�	�z�5ߋ��ߗ���PONITO�R�G ?kK  � 	EXEC�1o�2�3�4��5��@�7�8
�9o��� ��(��4��@��L� ��X��d��p��|⪂�2��2��2��2���2��2��2��2���2��2��3��3��3(�#AR_GRP_SV 1��[� (�1@2�����<�X���gs��`8Ͽ�v>RM�A_D�sҔN��ION_D�B-@�1Ml  �� �FH" �Zl �/� sFH~��N   5�c ��/]FI-u�d1}E���)P�L_NAME �!�E� �!D�efault P�ersonali�ty (from� FD)b (RR�2�� 1�L��XL�p�X  d�-?Qc u������� //)/;/M/_/q/�/�/�/EC2)�/�/�/ ??,?>?P?b?t?EB<�/�?�?�?�?�?�?�
OO.O@OROdO��6�?�N
�O�O�P�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_�O�O2oDoVoho zo�o�o�o�o�o�o�o 
.@o!ov� ���������*�<�N�`�r������ FR GT��G�M���  #�ÏՍ�d���� ���(�6������
� �m�~�h����� ������ğ֟������:���
�]�m����	`������į��:�oA������ A�  /���P����r��� ����^�˿ݿȿ��t%��R�� 1��	�X ��, �� ��� a� @D7�  t�?�z�`��?� |��A/��xt�{	��;�	l���	 �x7J������ ^�� �<�@����� ��·�K���K ��K=*��J���J���J9��
��ԏC߷�t�@{;S�\��(Ehє���.��I����ڌ���T;f��ґ�$��3���/�  �@���������$�  >����ӧU���x`���� �
����Ǌ��� �  {  @T�}����  �H ��l�ϊ�-�	'�� � ��I� �  �<��+�:�È��È�=�����0Ӂ���N �[��n �@���f����f��k���,�av�  '������@2��@�0@�Ш����C��Cb C���\C������Gs�@f �� I I����� )�Bb �$/�!��L�Dz �o�ߓ~��0���( �� -��������!9�D�  |9�恀?�ffG�*<� }�q�"1�89��>��bp$��(�(9��P��	�������>�?���9�x9�W�<
6�b<߈;܍��<�ê<���<�^��I/��A�{��fÌ�,��?fff?_�?&�� T�@�.�"��J<?�\��"N\�6���!��(�|� �/z��/j'��[0?? T???x?c?�?�?�?�?0�?�?6��%F���? 2O�?VO�/wO�)IO�O�EHG@ G@0~9�G�� G}� �O�O�O_	_B_-_f_�Q_BL9�B[�A w_[_�_b��_�[�_�� mO3o�OZo�_~o�o�o<�o���b��PV( @|po	lo-*cU�ߡA���r5�9�CP�Lo�}?����#��6���W9���6�Cv�q�CH3� j�t�����q�����|^(�hA� �ALf�fA]��?�$��?��;�°�u�æ�)�	�ff��C�#s�
���g\)�"��33C�
�����<�؎�G�B������L�B�s�����	";�H��ۚG��!G���WIYE���C�+�8��I۪I�5��HgMG�3�E��RC�j=�x�
�pI����G��fIV=�?E<YD�C<� ݟȟ����7�"�[� F��j�������ٯį ���!��E�0�i�T� f�����ÿ���ҿ� ���A�,�e�Pω�t� �Ϙ��ϼ������+� �O�:�s�^߃ߩߔ� �߸������ �9�$� 6�o�Z��~����� �������5� �Y�D� }�h����������������
C.(䁳3��/"���<���t��q3ǭ8����q4M�gu���q�Vw�Q�
4p�+4�]$$dR�Pv���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/�/X�/�/�/  %��/ �/+??O?:?s?/�_0�?�?�?�;�?�?@O�? OFO4O�rLO�^O�O�O�O�O�O�J � 2 Fs�wGwT�V�M�uaBO�|r�pp�C��S@�R_�poy_�_�_l�_o \!�W�Ƀh_oo(o�z?_���@@�z�D��p�pk1�p�~
 6o�o�o�o �o�o�o);M�_q�ڊsa �����D��$M�R_CABLE �2�� �]��T�LaMa?��PMaLb�p�Z���&P�C�p?aO4>ߔB���?aY�4?`?aE�h�\?f��v�l  ���&P�v�wdN��{0��$s8<ca��F�� 6��H�XT��6P?`C$��Č��n���	?`'z�"�,����� ��&P���C���=��������?`)z��~։��s9��T� ,�>���b�������Ɵ ��Ο3�.��P�(�:�@��^���j��#?`�� ����<h�H�Z�l��<h*��** ��sOM ��y����B�B�6-�%% 23456�78901ɿ۵ �ƿ���?`�?`AQ�?`?a
�z��not sent� ���W��TESTFECS7ALG� eg;jAQ�d��ga%�
���@��?d�r�̹�������� 9UD1�:\mainte�nances.x�mS�.�@�vj��DEFAULT��\�rGRP 2�^��  p?`�J�?e  �%1s�t mechan�ical che�ck�?a���������E��Z��(�:�L�^�?b��co�ntroller �Ԍ��߰��D���`�� ��$�s�M��L�?b"8b���v��B������������/�C}�a�6�����dv���s�C���ge��. battery�&��E	S(:L^pܿ	|�duiz�ab;let  D�а�R����/"/4/s��grgeas�>gf�r#!-?`|!�/�E��/��/�/�/�/s�
�oai,�g/y/�/�/@t?�?�?�?�?s��
$�?f�W��1<?`AO�E
c?8OJO\OnO��O�t��?O���'O�O_ _2_D_s�OverhauE�6�L��R x?`�Q�_���O�_�_�_�_o?`$�_0o����_o �_�o�o�o�o�oo �o?oQocoJ\n ���o�)� �"�4�F���|�� k��ď֏����[� 0�B���f��������� ��ҟ!���E�W�,�{� P�b�t�����矼�� ��A��(�:�L�^� ����ѯ㯸��ܿ�  ��$�s�Hϗ���~� Ϳ�ϴ�������9�� ]�o�Dߓ�h�zߌߞ� ������#�5�G���.� @�R�d�v��ߚ����� �������*�y��� `���O���������� ��?�&u�J��n �����); _4FXj|� ���%�// 0/B/�f/���/� �/�/�/�/?W/,?{/ �/b?�/�?�?�?�?�? ?�?A?S?(Ow?LO^O pO�O�O�?�OOO+O �O_$_6_H_Z_�O~_ �O�O�O�_�_�_�_o8 o�PeR	 T"oOo aoso�_�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
���  ��Q?� ; @eQ �oW� i�{�eVC�����̟bXw*�** �Q �V��� �2�D��h�8z��������_�S ������կ7�I� [�����ɯ/���ǿٿ #���!�3�}����� {ύϟ��s������� C�U�g��S�e�w�9�@�߭߿�	��eUeQ��$MR_HIS�T 2��U��� 
 \jR$ 2�34567890�1*�2����)�9 c_���R��a_���� �����=�O�a��*� x�����r����� ��9��]o&�J �����#� G�k}4�Z��SKCFMAP � �U�����Z��ONREL  �����лEXC/FENB'
���!FNC$/$JO�GOVLIM'd��m �KEY'zp%y%_PAN(��"�"�RUN`,�p%�SFSPD�TYPD(%�SI�GN/$T1MO�Tb/!�_CE_GRP 1��U�"�:`��n?Z [?�?�؆?�?~?�?�? �?!O�?EO�?:O{O2O �O�OhO�O�O�O_�O /_�O(_e__�_�_�_ �_v_�_�_�_o�׻QZ_EDIT4���#TCOM_C_FG 1��'%�to�o�o 
Ua_A�RC_!"��O)T�_MN_MODE�6�Lj_SPL��o2&UAP_CP�L�o3$NOCHE�CK ?� � Rdv� ���������*�<�N�`��NO_?WAIT_L 7Jg650NT]a���UzZ��_ERR?12���ф��	���-����R�d����`O�����| �O��
aC 	=�����?��y��0�¶��lW<� �� ?��j�ϟj����قPA�RAMႳ��N�
oQ�h�o��� = e���� ��گ�ȯ��"�4��0X�j�F�g蜿���A�ҿ�"ODRDS�P�c6/(OFFS?ET_CAR@`�o��DIS��S_�A�`ARK7KiO�PEN_FILE�4�1�aKf�`OPT?ION_IO�/�!���M_PRG %�%$*����h��WOT��E7�O����Z��  %��"�÷"�G	 �W"�Z����RG_DS�BL  ���ˊ���RIENTkTO ZC����A �U�`IM�_D���O��V~�LCT ����Gbԛa�Zd��_�PEX�`7�*�RA-T�g d/%*���UP ���{��������������/$PAL�������_POS_CHU��7����2>3�L��XL�p��$�ÿU�g�y��� ������������	 -?Qcu����Y2C���" 4FXj|�� ���� //$/6/@H/Z/l/~/�Y�� �.��/�/ςP�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO�/ �/LO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_)O;O�_�_�_�_�_ �_�_o o2oDoVoho�zo�o�o�_��� �o�m ���(�"{ BPw�m�m���~�jw8��w���� ��2�T��p��w���H��t	`���̏ޏ��:�o������ �2��pA�   I��j�`������ ���џ���@���#�)�Or�1����� 8�>��, �\Ԡ�~� @D�  ��?���~�?� ���!�D������%G� � ;�	l��	 ��x�J젌����� ��<� ��� ���2�H(��H�3k7HSM5G��22G���GN�3%�R��oR�d��2�Cf��a��{������������3��-¸��4��>����𚿬���3�A�q�½{q�!ª��ֱ� "�(«�p=�2����� ��_{  @�Њ��_�  ��Њ��2��ς�	'� �� ��I� ��  �V���=�������˖ß���  �y��n @"��]�<߭�"��������N�Д߇  '�Ь�w�ӰC>��C��\C߰���Ϲ��ߤ!���@%�4���/��2�~�B��B�I�;�)�j客z+���쿱����������( �� -��#�������!�]�9�|�  q�?�ffaH�Z��� ������"��8� ����>�|P$��}�(� ��P��������\�?���� x� ���<
6�b<߈;܍��<�ê<���<�^�*�gv�A)ۙ�脣��F��?fff?}�?&�� ��@�.���J<?�\��N\��)������� ����ޤy�N9 r]������ �/&/�J/5/n/��	g/�/c(G@� G@0i�G�� G}���/??<?�'?`?K?�?o?BL
i�B��A�?y?�?|� �?K�?ů�/QO�/xO��?�O�O�O�Om��bs��n�t @|�O '_�OK_6_H_�_�3��!A��RS�i�Cn_�_xj_0O�]?��o�oAo,où�Wi����ToC���`CH�Qo>Jd�`a�a@�Iܚ>(hA�� �ALffA�]��?�$�?����ź°u��æ�)�	ff���C�#�
ܢopg\)��3�3C�
������<��nG��B���L��B�s�����	0źH����G��!G���WIYE����C�+�½I�۪I�5�H�gMG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo�� �
��U�@�y�d��� ������я����� ?�*�c�N���r����� ���̟��)��9� _�J���n�����˯�� �گ�%��I�4�m� X���|���ǿ���ֿ ���3��W�B�Tύ� xϱϜ���������	� /��S�>�w�bߛ߆� �ߪ߼�������=��(�a�L�(q���)����Z�������a3�8�������a4Mgux�����a�VwQ��(�4p�+4�]B�B���p�����������UPbP���Q O%x�1[FjR�������  C���I 4mX�8
O������.//>/d/R/�Rj/|/�/�/�/�/�/:  2� Fs�gGT]�&6�M�eBmpX�R�P�aC��3@�_ p?�?�?�?�?�?�=�S�OO)O;OMO�c�?���@@�jJ��`�`�1�`�^
 TO�O�O �O�O�O_#_5_G_Y_�k_}_�_�_�j�A �����D��$�PARAM_ME�NU ?B���  �DEFPULS�E�[	WAIT�TMOUTkR�CVo SH�ELL_WRK.�$CUR_STY�L`DlOPT�Z1ZoPTBooibC�?oR_DECSN `���l�o�o�o &OJ\n������QSSREL_ID  >��
1��uUSE_P�ROG %�Z%8�@��sCCR` ��
1�SS�_HOST7 !�Z!X����M�T _���x�������L�_TIME�b �h��PGDE�BUG�p�[�sGI�NP_FLMSK��E�T� V�G�PG�Ar� 5��?��CyHS�D�TYPE�\�0��
�3�.� @�R�{�v�����ï�� Я����*�S�N� `�r����������޿ ��+�&�8�J�s�n���ϒϻ�G�WORD� ?	�[
 	�PR2��MA9I�`�SU�a��cTEԀ���	Sd�COL��C߸��L� C�~��h�d*�TRACE�CTL 1�B���Q ��m n'��0�ށ�_DT Q�B������D � ���q����
�����1�@� �@⨐�@�@�U � �	����U�������&�U�.�������U���&��.��6�U�>��F�
H�H�H����������K H� ������5��������U�������&��.��6��>�U�g��y���G�������Ѯ��� ���� ��������/�A�S� e�w��������������������O
��OO�Ug��X��XXX
X�Xf�����V�V�V�V���V��V��V��V���V��V��V���!�������@�� �� 2DNhz �f����-�?� ���?�?�?�������� ��d5(O:OLO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�P�$Or������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~�f���� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo��o�o�o�o�o�a�$�PGTRACEL�EN  �a  ���`���f_UP �/���q'pq� p�a_CFG7 �u	s�a p�LtLtfqw|pqz  �qu�4rDEFSPD ��?|�ap���`H_CONFI�G �us U�`�`d�t��b �a�qP�t�q���`��`IN7pT�RL �?}_q8l�u�PE�u��w�qLt�qqv�`WLID8s�?}	v��LLB 1��y� ��B�pB94Ńqv �އ�؏	�s << �a?��'�� �A�o�U�w������� ۟��ӟ��#�	�+�Y�v�񂍯����ï
���������/�u�GRoP 1ƪ��a�@�j��hs��aA�
D��� D@� Cŀ7 @�٭^�t�q0�����q�p���.� ���Ⱦ´���ʻB�)�	���?�)��c��a>��>��,��Ϻ��ζ� =49X=H�9�� 
����@�+�d�O����s߬�o߼�����  #Dz���`
��8� ��H�n�Y��}��� ����������4��X��C�|���)��
V�7.10beta�1Xv A������!�����?�!G�>\=�y�#��{33A!��@��͵���8wA��@_� A�s�@Ls���� ��"4FX�LsApLry�ā�_��@l�ͯ@�33q�`s���k��Anff��a��ھ��o)�x�� �a r�T�n�t�����	t�KNOW_M�  |uGvz�SV7 ��z�r� &����>/�/PG/�a��y�MM���{� ���	^u (l+/�/',_t�@XLs	����@���%�"�4�.N�z�MRM��|-TU�y�c?u;e�OADBANFW�D~x�STM�1 �1�y�4Garra_B�2Sem��?~s�;Co�2��O�7��3Antena�_Full @� �VODe�qH��^OpO �O�O�O�O�O�O!_ _ _W_6_H_�_l_~_�_��b�72�<�!4�_ � �<�_�_N�3 �_�_
oo�749oKo]ooo�75�o�o�o�o��76�o�o�77 2DVh�78��X���7MA�0���swwOVLD � �{�/a�2P�ARNUM  p�;]��u�SCH*� 8�
����ω�3�UPD��[�ܵ+�>wu_CMP_r -���0�'�5C�ER�_CHKQ���`�1�"e�N�`�RS>0��?G�_MO�?_���#u_RES_G
�0��{
Ϳ@�3� d�W���{�������� կ���*�����P��O��8`l��� ����`��ʿϿ��` �	���1p)�H�M� ��phχό���p��x�����V 1��5|�1�!@`y�ŒTHR_INR>0�/�Z"�5d:�MASmSG� Z[�MNF��y�MON_QUEUE ��5�6ӐV~  #tNH�U��qN�ֲ���END�����EXE������BE������OPT�IO������PROGRAM %���%��߰���TA�SK_I,�>�OCFG ά�]���^��DATAu#������! 2 ����R�d�0v�����:� ��� ������������ �2DV	�INFO
u#� ���Ԕ$�� ����
.@ Rdv�����@��/as x� �c ;���ȀK_������S&ENB�-�b-&q�&2�/�(G���2�b+ X,�		��=���/��@��P4$��0��99)�N'_E?DIT ���W?|i?��WERFL��-ӱ3RGADJ K�F:A@�5?Ӑ��5Wј6��]!֐���?�  Bz�WӐ<11�ҁ%�%O�8;��50!2Y��7�	H��l0��,�BP�0�s�@�0�M*�@=/�B **:�B�OH�F�O2��D��A�� �O�@O	_,X��%���H�q��O$_r_ 0_�_���Q@WA��>] �_�_�_o�_o�_�_ 
o�o.o�ojodovo�o �o�o�o�o�o\X B<N�r��� �4��0���&��� J������������� ����x�"�t�^�X� j�䟎���ʟğ֟P� ��L�6�0�B���f��� ������(�ү$��� ���>���z�t��� � �������l��h�R�L�^�DX	���ώ0x�� ���t$ :߀L��o�
ߓߥ��7P?REF ��:�0�
�5IORIT�YX�M6��1MPD�SPV�:n" �UT���C�6ODUCT���F:��NFOG[@_TG�0��J:�?�HIBIT_D�O�8��TOENT� 1�F; (!AF_INE*������!tcp|���!ud��~8�!icm'���N?�XY�3�F<��1)� �A�����0��������� ��' ]D�h�������*>��3��9n"OTfN�3>����B�G!/�LC��4�;LFJ�AB,  � ��F!//%/7/�5�F�Z�w/�/�/�/��3&ENHAN�CE �2FBA�H+d�?�%;��������Ӓ1�1POR_T_NUM+��0����1_CAR�TRE�@��q�S�KSTA*��SL�GS�������C�Unothing?�?OO����0TEMP ��N�"O�E�0_a_?seiban|߅O xߕO�O�O�O�O_�O '__K_6_H_�_l_�_ �_�_�_�_�_�_#oo Go2okoVo�ozo�o�o �o�o�o�o1U @e�v���� �����Q�<�u�>.IVERSI	�L���� dis�able'2*KSA�VE �N�	�2670H771|�h��!�/��9�:� 	^�4�ϐ�	���e��͟ߟ�����9�D�C-Å]_y� 1������ő����Ǻ�/URGE� B��r�WFϠ��-��9��W����l:WRU�P_DELAY ��=n�WR_HOT %��7��/�p��R_NORM�ALO�V�_�����S�EMI��������Q/SKIPo��97��xf�=�b�a�sυ�H� �ʹ��ø�������� &��J�\�n�4�Fߤ� �������߲���� � F�X�j�0��|���� �������0�B�T� �x�f���������ãRBTIF�5���CVTMOU�7v�5���DCRo�}�� �T��A�:CC�av�C�>�;P�>�[a:�_��H�� �cÄ���^��?�S�`?kϻ4�HϘ��� <
6b<�߈;܍�>�u.�>*��<��ǪP0���2DVhz��������,GR�DIO_TYPE�  v��/ED�� T_CFG ���-�BH]�E�P)�2��+ ��B�u �/�*��/ �?�/%?=�/V?� }?�Ϟ?���?�?�?�? �?O
O@O*Gl?qO�� 8O�O�O�O�O�O�O�O �O_<_^Oc_�O�__ �_�_�_�_�_o�_&o H_Mol_o�oo�o�o �o�o�o�o�o"DoI ho*j���� ���.3�E��f�  ���x��������ҏ �*�/�N��b�P��� t�����Ο��ޟ�:��+���R'INT 2��R��!�1G;�� i�{��"���8f�0 ��ӫ��� ���M�;�q�W��� ����˿���տ�%� �I�7�m��eϣϑ� �ϵ�������!��E� 3�i�{�aߟߍ��߱߀��������A���E�FPOS1 1�~!)  x� ��n#���������� ����/��S���w�� ��6�����l����� ��=O����6�� �V�z� 9 �]����R d���#/�G/� k//h/�/</�/`/�/ �/??�/�/?g?R? �?&?�?J?�?n?�?	O �?-O�?QO�?uO�O"O 4OnO�O�O�O�O_�O ;_�O8_q__�_0_�_ T_�_�_�_�_�_7o"o [o�_oo�o>o�o�o to�o�o!�oEW�o >���^�� ���A��e� ��� $�����Z�l����� +�ƏO��s��p��� D�͟h�񟌟�'� ԟ�o�Z���.���R� ۯv�د���5�ЯY� ��}���*�<�v�׿¿ ����Ϻ�C�޿@�y�<�e�2 1�q�� -�g�����	��-��� Q���N߇�"߫�F��� j��ߎߠ߲���M�8� q���0��T���� �����7���[���� �T�������t����� !��W��{� :�^p�� A�e �$�� Z�~/�+/�� �$/�/p/�/D/�/h/ �/�/�/'?�/K?�/o? 
?�?.?@?R?�?�?�? O�?5O�?YO�?VO�O *O�ONO�OrO�O�O�O �O�OU_@_y__�_8_ �_\_�_�_�_o�_?o �_co�_o"o\o�o�o �o|o�o)�o&_ �o��B�fx ��%��I��m�� ��,���Ǐb�돆�� ��3�Ώ���,���x� ��L�՟p�������/� ʟS��w�����ϓ�3 1��H�Z��� ���6�<�Z���~�� {���O�ؿs����� � ��Ϳ߿�z�eϞ�9� ��]��ρ���߷�@� ��d��ψ�#�5�G߁� ������*���N��� K����C���g��� ������J�5�n�	� ��-���Q������� ��4��X��Q ���q��� T�x�7� [m�//>/� b/��/!/�/�/W/�/ {/?�/(?�/�/�/!? �?m?�?A?�?e?�?�? �?$O�?HO�?lOO�O +O=OOO�O�O�O_�O 2_�OV_�OS_�_'_�_ K_�_o_�_�_�_�_�_ Ro=ovoo�o5o�oYo �o�o�o�o<�o` �oY���y ��&��#�\��������?�ȏ����4 1�˯u�����?�*� c�i���"���F���� |����)�ğM���� �F�����˯f�﯊� ����I��m���� ,���P�b�t������ 3�οW��{��xϱ� L���p��ϔ�߸��� ���w�bߛ�6߿�Z� ��~�����=���a� �߅� �2�D�~����� ���'���K���H��� ���@���d������� ����G2k�* �N����1 �U�N�� �n��/�/Q/ �u//�/4/�/X/j/ |/�/??;?�/_?�/ �??�?�?T?�?x?O �?%O�?�?�?OOjO �O>O�ObO�O�O�O!_ �OE_�Oi__�_(_:_ L_�_�_�_o�_/o�_ So�_Po�o$o�oHo�o�lo�oۏ�5 1� ���o�o�olW��o �O�s���2� �V��z��'�9�s� ԏ���������@�ۏ =�v����5���Y�� }�����۟<�'�`��� �����C���ޯy�� ��&���J����	�C� ����ȿc�쿇�ϫ� �F��j�ώ�)ϲ� M�_�qϫ����0��� T���x��u߮�I��� m��ߑ�������� t�_��3��W���{� �����:���^���� �/�A�{����� �� $��H��E~� =�a����� D/h�'�K ���
/�./�R/ ��/K/�/�/�/k/ �/�/?�/?N?�/r? ?�?1?�?U?g?y?�? O�?8O�?\O�?�OO }O�OQO�OuO�O�O"_<t6 1�%�O �O_�_�_�_�O�_|_ o�_o;o�__o�_�o o�oBoTofo�o�o %�oI�omj� >�b����� ��i�T���(���L� Տp�ҏ���/�ʏS� �w��$�6�p�џ�� �������=�؟:�s� ���2���V�߯z��� ��د9�$�]������ ��@���ۿv�����#� ��G�����@ϡό� ��`��τ�ߨ�
�C� ��g�ߋ�&߯�J�\� nߨ�	���-���Q��� u��r��F���j��� ����������q�\� ��0���T���x��� ��7��[��, >x����!� E�B{�:� ^�����A/,/ e/ /�/$/�/H/�/�/ ~/?�/+?�/O?5_GT7 1�R_�/?H? �?�?�?�/O�?2O�? /OhOO�O'O�OKO�O oO�O�O�O.__R_�O v__�_5_�_�_k_�_ �_o�_<o�_�_�_5o �o�o�oUo�oyo�o �o8�o\�o�� ?Qc���"�� F��j��g���;�ď _�菃������ˏ� f�Q���%���I�ҟm� ϟ���,�ǟP��t� �!�3�m�ί��򯍯 ���:�կ7�p���� /���S�ܿw�����տ 6�!�Z���~�Ϣ�=� ����s��ϗ� ߻�D� �����=ߞ߉���]� �߁�
���@���d� �߈�#��G�Y�k�� ���*���N���r�� o���C���g����� ������nY�- �Q�u��4��X�|b?t48 1�?);u�� /;/�_/�\/�/ 0/�/T/�/x/?�/�/ �/�/[?F???�?>? �?b?�?�?�?!O�?EO �?iOOO(ObO�O�O �O�O_�O/_�O,_e_  _�_$_�_H_�_l_~_ �_�_+ooOo�_soo �o2o�o�oho�o�o �o9�o�o�o2�~ �R�v���5� �Y��}����<�N� `���������C�ޏ g��d���8���\�� ��	�����ȟ�c�N� ��"���F�ϯj�̯� ��)�įM��q��� 0�j�˿��ￊ�Ϯ� 7�ҿ4�m�ϑ�,ϵ� P���tφϘ���3�� W���{�ߟ�:ߜ��� p��ߔ���A�����  �:����Z���~� ����=���a����� �����MASKW 1����������XNO  ����� MOTE �   N_C�FG �Y�����PL_RANG�UP���OWE/R ��� ��A��*SYST�EM*P�V9.3�044 �1/9�/2020 A� �g ���RE�START_T �  , $F�LAG� $DS�B_SIGNAL�� $UP_C�ND4P��RS2�32r � �$COMMEN�T $DEVICEUSE4�PEEC$PAR�ITY4OPBI�TS4FLOWC�ONTRO3TI�MEOUe6CUz�M4AUXT���5INTERFA�CsTATU�o �KCH� t $O�LD_yC_SW� 'FREEF?ROMSIZ ��ARGET_DI�R 	$UP?DT_MAP"� TSK_ENB"�EXP:*#!jF�AUL EV!�RV_DATA��  $n E��   	$VA�LU�! 	j&G�RP_  � {!A  2� �SCR�	� �$ITP�_�" $NU�M� OUP� �#T�OT_AX��#D�SP�&JOGLI��FINE_PC�d�OND�%$�UM�K5 _M�IR1!4PP TN�?8APL"G0_EXb0<$�!� 814�!{PGw6BRKH��;&NC� IS :�  �2TYP� �2��"P+ Ds�#;0B�SOC�&R N�5DUMMY164�"�SV_CODE_�OP�SFSPD__OVRD�2^�LDB3ORGT-P; LEFF�0<G�� OV5SFTJR3UNWC!SFpF5�%3UFRA�JTO~�LCHDLY7RECOVD'� �WS* �0�E0RO��10_p@  � @��S NVwERT"OFS�@9C� "FWD8A�D<4A�1ENABZ6�0�TR3$1_`1F�DO[6MB_CM��!FPB� BL_MP��!2hRnQ2xCV� "' } �#PBGiW|8AMz3\P��U�B�__M�P�M� �1�AOT$CA� �PD�2�PHBK+!:&a�IO�4 eIDX+bPPAj?a$i�Od7e�U7a�CDVC_DBG"�a;!&�`�B5�e1�j�S�ey3�f�@ATIO� ���AU�c� �S&�AB
0Y.#0 �D��X!� _�:&?SUBCPU%0SIN_RS�T, �1N|�S�T!�1$HW_C1�"]q.`<�v�Q$AT! � ��$UNIT�4|�p�pATTRI= ��r0CYCL3N�ECA�bL3FLT?R_2_FI9a7��c,!LP;CH�K_�SCT>3F�_�wF_�|8��zFqS+�R�rCHAGp��y��R�x�RSD��@'�1E#&7`_T��XPRO�`@S�E�MPER_0�3T�f�]p� f��P�D�IAG;%RAIL�AC�c4rM� LOh�0�A�65�"PS�"b�2 -`�e�SPR�`MS.  �W�Ctazf	�CFUNC�2��RINS_T�.!(�w��� S_� �0�P�� 	d���WARL0bCBL'CUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!2��8�3�TID�S���!� $CE_R�IA !5AFDpPbC~��@��T2 �1C9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@H�RDYOL1	PRG�8�H��>1(�ҥM�ULSE =#Sw3.��$JJJ6BKG�FKFAN_ALMsLV3R�WRNY��HARD�0+&_P� "��2Q���!�5_,�@:&AU�Rk��?TO_SBRvb���� ƺ�pvc�޳MPINF�@�q�)�N��REG'd~0V) x0R�C�1DAL_ �\2FL�u�2$M@Ԑ(�#S��P� `�6g�CMt`NF�qsCONIP�q5" �IP�P 9a3$Y��! �"�!�� �o3EaGP��#@��AR� ��c�52�����|5A�XE�'ROB�*R�ED�&WR�@�1_=��3SY�0ѥ0_�Si�WRI�@�ƅpST�#��0*@� B�q	���3��� B� ��A��3�D�POTOr�� �@ARY�#`��!��d�!1FI�0~�$LINK���GTH�B T_����A��6�"/�X�YZ+"9�7G�OFIF�@�.�"���	B� l����A3$ ��FI�p���4�4l��$_Jd�"(B �,a������8�"q�������Ck6D�UR��94�TURBT�XZ�N����Xx��P��FL/�@s���l�P��30�"Q W1� K
0M:$�53]q7�SuD�Sw#ORQɆ�!�����Q7��0O[�ND�=#8�!#�1OVE8��M���R��R�Q!P.!P! OAN}q	�R����990 � �brJ9V��Ø�v�!ER1��	B8�E�@n D�A��p�嘕Ă���v�AX�C�"��`�q �s���0~ 3�~F�~e�~�~E�~1��~Ҡ{Ҡ �Ҡ�Ҡ�Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�!�)DEBU}s$�x���삼!R*�AB��a8A2V`|r 
�"�c���%�Q7 �7�173�7F�7 e�7�7E����\���LAB����yp�cGRO�p��}��PB_ҁ ��̓ ��ð�6�1���5���6AND��8p�a3���-G �Q����AH0�PH�p2�NTd��Cs@VEL؁�}A�~�F�SERVEs@N�� $����A!�!�@POR}�KP��иA���@���	�  $�BTREQ�
�CH��@
�GƄ�2	�Eb��_ � lb��Q�ERR��RI�P�@�NFQTOQ�� L�P}��YVĀG�E%�\��CRE� � ,�A�EP
��RA�Q 23 d�R7c�T�@7 ��$F ׂ4��m �DOC��P�  8[CO�UNT���@��FZ�N_CFG�A 4�p%��rT\zs�a��#`pJp c%d�� �� MGp+����`0�OGp�eFAq����cX8еk�ioQ�¤'ѴDp8�Pz����SHELA�-b� 5��B_wBAS\RSR$Ɗ`�2�S��L�!p1T�W!p2Dz3Dz4DzU5Dz6Dz7Dz8�WqROO���P�1�3NL�� �AB�C
�n"pACK�&IN�P	T+�W�U��	�k��y�_PU8�~�|�OU�CP��%�s�Vl����YTPFWD_KcARKQ-�:PRE�D��P����QUE�$�Ā9 )���~���I U��#s/���@�/�SEM1ǆ1�An�aSTY�tSO����DI�q��Qc��X_TM9�MANsRQ �/�END���$KEYSWI�TCH2�G����H}E)�BEATMz�PE��LEJR���0Jx�UF�F��G�S��DO_HOM��Olz��pEFPR��PSbJі��uC��O��<7P�QOV_M��}�c�IOCM���1���QsHK��# D,�&�a`U2R���M��a�r +�FORC*�WAR�hbs�OM��  @��$�㰰U��P�1���g���3��4��E��S�POW�Lz�<�R%�UNLO�0T��ED��  ��SNP��S.b; 0N�ADDa`z��$SIZ*�$�VA�0�UMULTCIP�r�P���Az� � $���ƒ���SQc�1C<FPv�FRIFr�PaSw���ʔf�NF#�ODBUx�R@w���0���F��:�IAh��Ƙ�������S"p��� �  �cRTE����SGL.�T�x�&C`Gõ3a�/�OSTMT��`�P����BW9 0�SHO�Wh�qBANt�TPo���E�������@V_Gsb �$PC�0�PokFBv�P��SP���A�p����D��rb�� �+QA002D.ҝ�6ק�6ױ��6׻�6�54�64�7�4�84�94�A4�B�4و�6ׇ17�}�6�F 4� ��@�����Z��T��t�1��1��1��U1��1��1��1��U1��1��1��23�U2@�2M�2Z�2g�U2t�2��2��2��U2��2��2��2��U2��2��2��33٨���M�3Z�3g�3�t�3��3��3��3���3��3��3��3���3��3��43�4�@�4M�4Z�4g�4�t�4��4��4��4���4��4��4��4���4��4��53�5�@�5M�5Z�5g�5�t�5��5��5��5���5��5��5��5���5��5��63�6�@�6M�6Z�6g�6�t�6��6��6��6���6��6��6��6���6��6��73�7�@�7M�7Z�7g�7�t�7��7��7��7���7��7��7��7���7��7�����Pzv�U�B �@ĳ09r
�����A �x �0R���  �BM�@RP�`�4Q_�PR�@[U�AR�J�DSMC��E2F�_U��=AhbYSL|�P�@ �  � ֲ>g�������iD��VALU>e�pL��A�HFZAID_L����EHI�JIh�$FILE_ ��D�dk$ǓVESA�Q� h�0!PE_BLCKz�.RI�7XD_CPUGY!�GY��Ic�O
TUB���R�  � PaW`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q��TJ��U�Q�T�Q�UH���T`�T�����T2L�_LIz��  �pG_O�T�P_EDI�U��T2�`7c �?bة�pBQh���]`B{C2 �! �%�`>��P��a�7aFTτ\�d݃TDC�PA��N`�`M�0�f�a�gT�H��U��d�3�gRx�q�9�ERVEЃt݃t	��a�p�`� "X -$EqLENЃRt݃Ep��pRAv��Y@W_�AtS1Eq�D2�wMIO?Q�S���pI��.B�A�y�4Ep�{DE<�u��LACE �C�CC�.B��_MA���v��w�TCV�:��wT,�;�Z�P�@��s�~��s�J�%A�M����J��R�uā�uQq2ѐ`���݁�s�JK��VK������	����J����JJ�JJ�AAL�<���<�6��:�5�cm�NA1a�m�,��DL�pa_\�Űѐ�aCF
��# `�0GROUP�@J�Բ��N�`C^�~ȐREQUIRr�ÀEBUu�Aq��$T�p2"��Bp�8�a	��d$ \?@qhoAPPR��CLB�
$H`N;�CLOD}`K�S�e`��u
�a.I�% �3�M�`�8l��_MG񱥠�C �"P����&���B{RK��NOLD����RTMO6a�ޭ��J6`�P>��p���p��pZ��pc��p6+�7+�<��QAq�d&� �lr���������PATH ��������qx�����9%0A��SCAub��l<���INDrUC�p��q�C�UM�Y�psP����A q/��/�E�/�PAYL�OA�J2L�0R'_AN�ap�L�Pz��v�jɆ���R_F2�LSHRt��LO�{�R�������ACRL_�q�����b�r�H�@B$H��^"�FLEX>�.`;BJ�f' P(��o��o+�p�aJDu( :Qcv�p�׀��f��po��|F1���-������]�E��*�<� N�`�r�����4�Q��� ����A�c���ɏۏ���T��2�X:A��� ���������)� ;�?�H�6�Z�c�u���t����J��) ��``��˟ݟ�`�0ATF�𑢀EL���a���J�(��JE۠C3TR��A�TN�1��HAND_VB�B>ѯ@�* $���F2���d�CS�W��<҉�+� $$M�����0ˡ�@ڡ������A�@ g����A)��A���@
˪A٫A� ��`P�˪D٫D�PȰG�P�)STͧ�!ک�!N�DY�P9���� #%��Fp���Ѫ���i� ���������P3�<��E�N�W�`�i�r�TP���, ��ԓ�� n�5m��1AS�YMص.@�ض+A������_`��	� ��D�&�8�J�\�n�Ju�&��ʧC�I��.S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R�� &T��3TWV�͢���&��ߪU��/�7Ӝ�f�0HR`ta-���QQ�1�DI��O��T����Q��. ; *"IAA*���$a`G�2C2cJ�$�H���P / � �ME�� Mb�R4AT�PPT�@� ��ua����P�l@zh�a�iT�@�� $�DUMMY1E�o$PS_D�RF��  ���f3�FL�A��YP���b}c?$GLB_T��U�uu`1�y���EQa0c X(���ST�����SBR�PM2�1_V��T$SV_ER��O_@KscsSCLpKrA��O'b��PGL�@EW��1s 4��a$Y,�Z,W�s怯��A�N`©�qU�u2 ���N�p�@$G�IU}$�q �14�s�p��3 qL���v^B}$F^B�E�vNEAR��N�K�F8���TANC�K��JOG��� �4��$JOI�NT��	a�qMS�ET��5  �wE�H�� S�J`�� ���6�  MU���?���LOCK�_FO����PBG�LVHGL�TE�ST_XM>���EMPt����r̀�$U�Гr��22���s,�3���Ҁ,��1MqCE���sM� �$KAR��M�ST�PDRA�pj�a�VcEC��{�e�IU,��41�HEԀTOOiL㠓V�RE��'IS3����6N�A�ACH���5��O��}c�d3���pS�I.�  @$R�AIL_BOXEz��ppROBO���?�pqHOWWA�R*���`�ROLM�bB���S��
��5�0O_F� !>ppHTML5�Q����"r�pڑ��]7m��R��O�ҡ8���v�z��vO�U��9 tpp(�1`4A�̀��PO֡]%PIP��N�����
�ڑS�,�����CORDEDҀް̠&5�XT��q) �� �O4` : D pOBP!"Ҁ{��j��cpj�^@$SYSj�ADR#�Pu`�TCH� ; M,��EN�RZ�Aف�_�t״�>����PVWVAPa<� � p��r�UP�REV_RT]1�$EDIT�VSHWR�7v;���J�q�@D_`#R�~+$HEADoAh�Pl�A$�KE�q��`CPSPD��J�MP��L�UV�TR��d=r�O�϶�I�S#CiNEx��$_TICK�b�AMX�b��HN-q> @t�������_GP��[�STYYѲ�LOqHb���Ҩ�?�
�G�ݵ%$���t=7pS !$Q��da�e�!`�fP�0�SQU�d� ��b�ATERC�y`Y��TS�@ �pCp����d�ė�%Oz`mcO�IZh�d�q�e�aPRM�0�a8����PUQH�g_DO=�ְXS���K�VAXIg�f�1�UR� ��$#��ȕ��� _����ET���Pۂ���5f�Fd�7g�A�!�1�d�9�2;����R|Al�о�� �#��5��#��#� )#�)i�>'i�N'i� ^&{����){����2��	C����C��WOiO{O܍D�qSSCp 7B hppDS(�k�f�`SP`�ATL ��I���¼bAD�DRES��B'�S�HIF��"�_2C�H#��I&p���TU&pI� C>��CUSTO��qV��IbDȲT,��0
�
��V塜X�R`E \����� f�7��tC�#	����F��irt�TX_SCREEl�F�P=��TINA�s�p���t  ��Q9_��0G T��fp ,⧱eqBp&uᦲu�$#�RRO'0R���p}�!���`�UE��GH ��0���`S�qN��RSM�k�UV�0���V~!�PS_�s�&@C�!�)�'C��Cǂ�z"� 2G�U�E�4Ibvr�&8�G+MTjPLDQ��Rp����
 �BBL�_�W�`R`J ��f�>2O�qJ2LE��U3"�T4RIG�H^3BRDxt�C'KGR�`�5TW��7>�1WIDTH�H�������a���U�Iu�EY��QaK Ad�p��A�J�
�4�BACKH��b�5|q�X`FOD�GLA-BS�?(X`I�˂�$UR(�9@�!I�_^`H4! L 	8�QR�_k��\B_`R�p͂����a�pIA)O�R`M��w0�Uj0�CRۂM�LUqM�C��� ERV�R�CP<��4NV`���GE=B#���]�t�LIP�E��E��Z)W@j'Xz'XԐ&Y5$[6$[7$[8	R���3�<���fԑŁSv��M�1USR�tOO <��^`U�r��rFO
�rPR�I��m����PTR�IP�m�UN[DO��P�p�� `m�4�l��0$����� QWB�P7�G �s�Tf�H�RbO	S�agfR��:">c��.qR��s�~�b*�~�#�UQ.qS�o�o�#8R)�>cOFF���p�T� �cOp �1R�t/tS�GU��P.q��JsETwn�1SUB*� f�_E_EXE��V��v>cWO>� U�`^g��WA'��P�q�!@� V_DB8�s�p�2SRT�`
�aV�Q�r��OR�N�uRAU��tT��ͷ�q_���W |�%�͸OWNA`޴�$SRCE � ��Dx��\��MPFIA�p��ESPD��� ���C���Gƒ�r-�5���!X `�`�r޴���COP�a$*�C`_w�������rCT�3�q���qƒp����@� Y"?SHADOW�ઓ~@�_UNSCA��8@��4M�DGDߑ��OEGAC�,Me��G�Z (0N�O�@�D<�PE�Bf��VW씸�RG���![ � ��VqEE#�aڒANG�$���c薴cڒLIM_X�c��c� �����#��`� ��bVyF� �s�VCCj�j��\ՒC{�RAl�p����RpNFA�i�%�E��Z`�G� ^0[�C`DqEĒ��� STEQ1 ���@�ꁻ@I��`+0�����`����P_�A6�r���K��!]�� 1Ҡ��� ��\��сCPC�@]�GDRIܐ\�͑V#�耴��D�TMY_UBY�T���c��F!����Y�븲���P�_V�y��LN�BMvQ1$��DEY��cEX�e��MU��5X�M� US�����P_R��b�P� ߖ=G��PACIr�ʐ f�ᔟ��c�´c���#B�EqB��aWrB�����^ ܀GBΐP����0C�R~`�`�_�0�@3!�1zr	4�e�R�SW��p��Yp��S�6�O�Q�1Ah� X�#�E�UE���Yp�`C�HKJ�`�@p���U� �EAN�ٖp�pXն��C�MRCV�!a U��@O��M�pC��	��s����REF *7
��������/��P ��@���@��b��֗�_Y��ژ��ۣ��Q$�3�����?��$b �����%���Q��$GROU� �c������ʠ]��I2^`0��U` 0_��I,�o � ULա`2��C&�rAaB�?�NT���������A���Q��K�L����õ���A���Q��T a$c� t�`MD�p8�H�U���SA�CMPE F  _�Rr�p@����9XS	��VGF/�b#_d, &�@M�P^0۰UF_C !���z �ROh0"+��p�@���0C�UREB����RI��
IN �p�����d��d�,�ca�INE�H�y��0V�a-�걗�3�W�������C��i�LO�}�z�@0�!�QNSI��݁����c$&�c$&.�X_PuE-YW+Z_M�ڒW�I�$�" �+�R�'rRSLre� �/�M
`�RE�C7�Gd�۰�� �ҭ�q����u��� �������S_P�V�nP�@�VIA�vf� �~pHDR�p�pJO�P��_$Z_UP��a_LOW�5�1J�dA���LINubEP�?�tc_i�1�1���@��G1@*�V�xg{ 5X�PATHP= X�CACH$��]E��yI�A��{�C�)�ID3FA�ETD��H��$HO�pO�b@�{�d6�F����<��p�PAGE�䁀�VP�°�(R_SI	Z��2TZ3�-X�0U̲q�MPRZ��IM5G���AD�Y��MRE��R7WGP���8�p��ASYN�BUF�VRTD��U�T7Q�LE_2�D-��U��`CҡU�1��Qu��UECCU��VEM��]EDb�GVIRC�Q�U�S��B�Q�LA��p�N�FOUN_�DIAuG�YRE�XYZ�cE�WѴh8�dpq2a`T��2�IM�a�V�|be��EGRABBr��Y�a�LERj��C4���FC-A�6504x��7u���2W����h'�`�CKLA�S_@l�BA��N@i I G��T��� @ݲ�մ$BAƠwj � !q�eb��uTYSp�H����2��I�t:b�f:��B)�EVE�����PK���fx��GI��pNO��2���#�H�O����k � @���
8�Pi�S�0�ޗ��RO�ACC�EL?0=���VR_�U7@�`��2�p��AR��PA��̎K�}D��REM_But7 T�rJMX ��l�t�$SSC��Uk[s�0G�QN@m� � �S�P�N�S��LEX�vn =T�ENAB 2¼W@��FLDRߨF�I�P�t�ߨ(Ğ����P2HFo� ���V
Q MV_PI��8T@�H���F@�Z� +�#��8�8#��sGAB���LOO󣎔�JCBx��w"SC�ON(P�PLANۀ�Dp�3F�d�v�9PէM��Q ;����SM0E�ɥ�8ɥWb 72$`<�8T��,`�RKh"ǁVANC�����R_Ou N@p (�-#<#c��c.2��w�A/�N@q 4������`	��^����w�N@r �hn���1^�&OF	F`|�p�`��`�D�EA�
�P,`SK��DMP6VIE��2�q w��@���rs < {���4����r{7��D���^L�CUST�U���t $G�TIT>1$PR\���OPTap ��VS)F�йsu�p�0`r�&� �0SMO"wvI�|�ĄJ����K�eQ_WB��wI����� @O3�@�X�VRxxmr��T����ZABC��y op�����)�
t�ZD$�CS;CH��z Lu��� �`�2�%PC ��7P�GN ��<��A��_�FUNH��@��ZI�Pw{I��LV�,SL��~�C��Z/MPCF��|��E�����X�DMY_L�NH�=�
D�� ��} $�A� ]�CMCM� C,SC�&!��P�� '$J���DQ��@�����������_�Q�,2����UX�a\�UXEUL��a�������(�:�(�J���F�TFL��w��Z�~�0+�6����Y@Dp � 8 $R�PU<��> EIGH����#?(�iֱ�b���et� �a����У$B�0�0@�	�_�SHIFD3-�RV2V`F�@��	$5��C�0��&!�������b
�sx�uD�T�R��V̱_��SsPH���!� ,���������4A�R;YP��%����%� �  �%!  *�H�(UN0�� �"�2�����K��q0GSPDak����P� �O����0��Ѱ��"!NGV�ER`q i�w+I_AIR�PURGE  i  i/�F`E�Tb� �+1h2ISOLC  �,��"� � �!��%��P+�_/*OBZ��Dm�?@�!�H771  34n?�?�9� `�E/#�)x� S23�2�� 1i�� LTEk@ PENDA�341l 1D3<*?� Maint�enance C�ons B�? F"�O,DNo UseMJOOnO�O�O�O8�O2�2NPO;/"j 19%�1CH=�8ɐ�.P		9Q_?!UD1:___�RSMAVAIL�/�/%�A!SR  �+��H�_�P�1�TVAL.&����P(.�YVL�}� �2i�� D?�P 	�/_oUQ No�orci�o�g�o�o �o�o�o*,> tb������ ���:�(�^�L��� p�������܏ʏ �� $��H�6�X�~�l��� ��Ɵ���؟����� D�2�h�V���z����� ���ԯ
���.��R� @�b�d�v�����п�� �����(�N�<�r��i�$SAF_D?O_PULS. j0Qp����CA� ��/%�&0SCR ��`�X�
�`�`
	14�1IAIE���b vo$�6� H�Z�l�~�ߢߴ��߰�������HS"��2%�����d1�(��8�rb��� @��"k�}���T�h� �J`���_ @��T7 �����#�~0�T D��0� Y�k�}����������� ����1CUg�y�O�Ef�p����  �5�;�o�� 1p��U�
�t���Di�������
  � ��*������ gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O7O<A���`OrO�O�O �O�O�O�O�O?O�_ ._@_R_d_v_�_�_�_�_�Q _�R0MJ To!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏJO��'�9�K� ]�o�������_ɟ۟ ����#�5�G�Y��_ �U�_�ҙ�����ϯ� ���)�;�M�_�m� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�;�?� q߮����������� ,�>�P�b�t�������������������Y��	�1234567�81h!B�!����F��� ��������������  ��;M_q ������� %7I[l*� ������// 1/C/U/g/y/�/�/�/ n��/�/	??-??? Q?c?u?�?�?�?�?�? �?�?O�/)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_O_ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �op_�o�o�o/ ASew���� �����o+�=�O� a�s���������͏ߏ ���'�9�K�]�� ��������ɟ۟��� �#�5�G�Y�k�}����������s�կ��w���0�L�CH�  Bpw�   ��=�2�� �} =�
~���  	�o�@ί��ǿٿ���r������@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖ�%� ����������&�8� J�\�n��������������"�Q�*�(����;�<M���D�~��  �]��w�*�Z򛱛�t C d�����*�`*���$SCR_GR�P 1*P�3� � }�*� 6��	 �
��<�+�*�'UC|@�Y�y�yD� W��!�y�	M-�10iA/7L �12345678k90��� 8���MT� � �
��	L��	Č� N
���Y���Dy�
M_	P������ ,���H�
 � ��1/@A/g/y/H���!T/�/P/�/3��+\���/B�S��,?�*2C4&Ad�R?  a@0j5N?�7?��7�&2R��?}:&F@ F�`�2�?�/�? �?OO-OSO>OwObO �O=j1�2�O�O�O�O�DB��O�O;_&___ J_�_n_�_�_�_�_�_ o�_%o�5j�eSgxo6���uo�o�b�1�B�|3�oh0�4j96j9B� w�$0Y̯@HtA�Nhcu$�/�%pp�drsqA ����z�q�x�� �� (&� *�2�D�V�oz�e��������ECLVL ; ����iqp�Q@��L_DEF�AULT �����փH�OTSTR�qq���MIPOWER�F��H���WF�DO� �RVENT 1Ɂ�Ɂ� L!D?UM_EIP������j!AF_I�NE‧���!FIT}�֞����!-/�� ��F�!�RPC_MAIN�G�)��5���Y�VI�Sb�t����ޯ!�TPѠPUկ��d�ͯ*�!
PMON?_PROXY+���Ae�v��D���fe��¿!RDM_S�RVÿ��g���!#R,*ϑ�h��Z�K!
[�M����iI����!RLSYN�C����8����!�ROS|���4���>�!
CE�MOTCOM?ߓ�k-����!	S�CONSd�ߒ�ly���!SҟWASRCݿ��m���"�!S�USB�#n�n�!S#TMC��o]�� ���ѳ����,����P�V�ICE_KL� ?%d� (%�SVCPRG1S�����2�������oD����4������5D��6;@��7c h�����9����%������� ��0����X��� ��-���U���} ��� /���H/�� �p/���/��F�/ ��n�/��?�� 8?���`?��/�?�� 6/�?��^/�?��/X� j��q���#OhO��lO �O{O�O�O�O�O�O�O  _2__V_A_z_e_�_ �_�_�_�_�_�_oo @o+odoOo�o�o�o�o �o�o�o�o*< `K�o���� ���&��J�5�n� Y���}���ȏ���^�_DEV d���MC:�4����GRP �2d���bx� 	� 
 ,V�ȡ�s�Z����� �������ߟ�� @�'�9�v�]�������@Я����۫Y����ܯI�1�4�]��� j�����˿F�Ŀ�� %�7��[�B��f�x� ���!���A����ۿ D�+�h�Oߌ�s߅��� ������
���@�'�d�v��	y��^��� ��������%��I�0� Y��f�����8����� ������3��T7]�e�����)� �
�.@�dK �o��!�9���!/G/���R/ �/�/�/�/�/"�/�/ ??C?*?<?y?`?�? ��?�?�?�?�?�?-O OQO8OaO�OnO�O�O �O�O�O_�O)_;_"_ __�?�_�_L_�_�_�_ �_�_o�_7oo0omo To�oxo�o�o�o�o�o !x_E�oU{b �������� /��S�:�w�^�p������я�d �XƿZI6 r���@Z��0�+�A����d�BjBA�=��������B����AZ.�A����+�A.��Q�B�����5\��i6�A��u��'��ǎ%�Ꮛ�%�PEGA_BAR�RA_ESTEI�RA����X�T����?=��=�X��7
�?��>�A����?������&����������AxP��f���U�'A�j���´�B��:�<�3�����jB]+a��T��%�T�腯d�ʐ���>�p�c?��7�Գ�T@6��A�_���0n�����·�Ak���۸I�K9�FA�G�����B!v,�-���C3�����pBM�>�#�b��(�Y�������HX��?L!���Q��B���AJߤ�Xk�@f�D3��O�A���������Yw���.B��B�;��C�H�z�B�?���6���-Ϙ������n��=]����V@����?,����Ö� վ���eAk�������OY�A��ㇾ��AB��J�;%�C$�4�aƿBXZ�9���
���ߘ��~��� �ԭ(��?^_��-\¯ԡ���گ���+������������ߔ�mᢧ��*נ�6�C>�ԯb���z���
��BM����s��x�U<~�߯7@6|=��C��$�6��� N�@���b�G���L��}������x7���~K@����V�+A>r�rF���������Y@+�@��<B��|�A��F����B)���,o�?ɇ���~0��0~�6�Z� Q������������Aߍ�]ܖ�A����ܺ����2[�����>�ȥA���=�³�NB ��$�w?�d�j��to�7\��
�.�%��Z�����A������*�@Ve��B� ������YN�#���BD�	����9A����gB#
q��3��C4#���,?[BVM����COLO�CA_PRENS�����&//J/ 8/n/\/~/�/�/ �/�/�/ ??D?2?T? �/�/�?�/z?�?�?�? �?O
O@O�?gO�?0O �O,O�O�O�O�O�O_ ZO?_~O_r_`_�_�_ �_�_�_�_2_oV_�_ Jo8ono\o�o�o�o�o 
o�o.o�o"F4 jX��o��~� z���B�0�f�� ���V�����Џҏ� ��>���e���.��� ������̟Ο���X� =�|��p�^������� ��ȯ�D��T��H� 6�l�Z���~�����ۿ ���Ϡ��D�2�h� Vό�ο���|����� 
����@�.�dߦϋ� ��T߾߬�������� �<�~�c��,��� ��������D�)�;� �����\��������� ���@���4"D FX�|���� ��0@BT ����z��/ �,//</���/� b/�/�/�/�/?�/(? j/O?�/?�??�?�? �?�?�? OB?'Of?�? ZOHO~OlO�O�O�O�O O�O>O�O2_ _V_D_ z_h_�_�_�O�__�_ 
o�_.ooRo@ovo�_ �o�ofo�obo�o�o *N�ou�o>� ������&�h M�����n������� ��ȏ��@�%�d��X� F�|�j��������,� ��<�֟0��T�B�x� f���ޟï������� �,��P�>�t����� گd�ο�����(� �Lώ�sϲ�<Ϧϔ� �ϸ�������$�f�K� ���~�lߢߐ��ߴ� ��,��#�������D� z�h��������(� ���
�,�.�@�v�d� ������ ������� (*<r����� b����$ z�q�J��� ���/R7/v / j/�z/�/�/�/�/�/ */?N/�/B?0?f?T? v?�?�?�??�?&?�? OO>O,ObOPOrO�O �?�O�?�O�O�O__ :_(_^_�O�_�_N_p_ J_�_�_�_o o6ox_ ]o�_&o�o~o�o�o�o �o�oPo5to�oh V�z����( �L�@�.�d�R��� v������$���� �<�*�`�N���Ə�� �t�ޟp����8� &�\�����L����� گȯ����4�v�[� ��$���|�����ֿĿ ��N�3�r���f�T� ��xϮϜ������� ���Ͼ�,�b�P߆�t� ������ߚ����� �(�^�L���ߩ��� r����� �����$� Z������J������� ������b���Y�� 2�z����� :^�R�b� v����6� *//N/</^/�/r/�/ ��//�/?�/&?? J?8?Z?�?�/�?�/p? �?�?�?�?"OOFO�? mOO6OXO2O�O�O�O �O�O_`OE_�O_x_ f_�_�_�_�_�_�_8_ o\_�_Po>otobo�o �o�o�oo�o4o�o( L:p^��o�o �� ��$��H� 6�l�����\�ƏX� ֏��� ��D���k� ��4�������ҟ�� ��^�C����v�d� ��������ί��6�� Z��N�<�r�`����� �����󿪿̿��� J�8�n�\ϒ�Կ���� �����������F�4� j߬ϑ���Z��߲��� �������B��i�� 2������������ J�p�A����t�b��� ��������"�F��� :��Jp^��� ���� 6$ FlZ����� ��/�2/ /B/h/ ��/�X/�/�/�/�/ 
?�/.?p/U?g??@? ?�?�?�?�?�?OH? -Ol?�?`ONOpOrO�O �O�O�O O_DO�O8_ &_\_J_l_n_�_�_�O �__�_o�_4o"oXo Foho�_�_�o�_�o�o �o�o0T�o{ �oD�@���� �,�nS�����t� ��������Ώ�F�+� j��^�L���p����� ��ܟ��B�̟6�$� Z�H�~�l����ɯۯ ��������2� �V�D��z��������$�SERV_MAI�L  ������ʴOUTPUT�ո�@�ʴRV 2j� � � (r�������=�ʴSAV�E���TOP10� 2� d 6 rƱ���� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t������n�YPY��F�ZN_CFG f��=���J���GRP 2���g� ,B  � A =�D;� �B �  B4~=�RB21I�oHELL��f�e�)�*�=�����%RSR��� ���&J5 G�k�������.�  ���/>/P/"\/ b�X/z"{ �U'
&"2�dh,g-�"E�HK 1S �/�/�/�/#?L?G? Y?k?�?�?�?�?�?�?��?�?$OO1OCO?OMM S�OD�FTOV_ENB�մ�e��"OW_R�EG_UI�O�IMIOFWDL~@��N�BWAIT��B�)��V��F��YTIM�E���G_VA԰_�A_�UNIT�C~Ve�L]C�@TRY�Ge��ʰMON_AL�IAS ?e�I%�he��oo&o8o Fj�_io{o�o�oJo�o �o�o�o�o/AS ew"����� ���+�=��N�s� ������T�͏ߏ�� ���9�K�]�o���,� ����ɟ۟ퟘ��#� 5�G��k�}������� ^�ׯ�����ʯC� U�g�y���6�����ӿ 忐����-�?�Q��� uχϙϫϽ�h����� ��)���M�_�q߃� ��@߹������ߚ�� %�7�I�[����� ����r������!�3� ��W�i�{���8����� ��������/AS e�����| �+=�as ��B����/ �'/9/K/]/o//�/ �/�/�/�/�/�/?#? 5?�/F?k?}?�?�?L? �?�?�?�?O�?1OCO UOgOyO$O�O�O�O�O �O�O	__-_?_�Oc_ u_�_�_�_V_�_�_�_�ooc�$SMO�N_DEFPRO�G &����Aa &�*SYSTEM*�obg $JO�0dRECALL �?}Ai ( ��}-copy m�db:*.* v�irt:\tmp�back\=>1�0.109.3.�21:9228 ��f:8664  ��`�o�o	t}1x�bfr:\�o'p�oA �o`r�r2ua%7�cP����q6ts:ord�erfil.dat�o�m�e�w�
��o 7��oR������ >Џa�s����)�;���ߟ���
xy�zrate 11 ����̟]�o�����=��:picku�p_barra_�esteira.�tp��emp��8�Z�����;����torno����ٯj��|��4�lace�1�C�ǁR����� �}:�sumir +�����ؿi�{����>��prens��H� Z������������K����j�|��<�furad��<�R�[�����ߑ�#�sem_recep1���H���0k�}�ߢ�co-�?�p������� }�61�� ����]�o����1 H�:�L��� ���&�����	m �$���H�U�� ��������dv� �.�D�Q��/�� ��O��f/x/�� �=/S/�/�/?�/ ?�/b?t?�?�,/9? O?�?�?O/�?�?M/ ^OpO�O�'�?K?�O �O _����I�Ol_ ~_�/�/,?�OY_�_�_ ?!?�_E?�_hozo�? �?2O�?Uo�o�oOO �oAO�odv��_�_ 6oQ���o�=o �`�r����o*<�o ޏ�������K\� n�����.��[�� ���#���G�ٟj�|�����$SNPX_�ASG 2�������o  0��%����Я  ?���PA�RAM ����� �	��P�ӤX�Ө$�������OFT_K�B_CFG  �ӣ����OPIN_�SIM  ����}���������R�VNORDY_DOO  )�U����QSTP_DSB�i��ϐ�SR ��� � &�#�D�O�O�:�TO�P_ON_ERR�ʿ��o�PTN ������A���RING_PR�My�ܲVCNT_�GP 2��!���x 	����X��ϰ#��Gߔ�VD��ROP 1��"�8� ��*߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�}�z��� ������������
 C@Rdv��� ���	*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?[?X?j?|? �?�?�?�?�?�?�?!O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo sopo�o�o�o�o�o�o �o 96HZl ~��������� �2�D�V�`�PRG_COUNTJ�s��{�ENB���}�M��L���_UP�D 1'�T  
k�����"�K� F�X�j���������۟ ֟���#��0�B�k� f�x���������ү�� ����C�>�P�b��� ������ӿο��� �(�:�c�^�pςϫ� �ϸ������� ��;� 6�H�Z߃�~ߐߢ��� �������� �2�[� V�h�z�������� ����
�3�.�@�R�{� v������������� *SN`r����t�_INFO� 1�Ҁ� 	 ���3�>�?�?� ?!�9 �C 	=����?��h���'�¶�l�>?�� A���@[� >�@� ?� A�@a �?���C�8�D��w�3������B� ���YSDEBUG������ dՉ�SP�_PASS��B�?+LOG ���� �  �a�  �сf!?UD1:\;$�<"_MPCA-셽/$�/�x!�/ 쁝&?SAV D)���%d!|"�%�(S�V�+TEM_TI_ME 1D'��W 0��쏄Ż
��',5M7MEMBOK  �сd �d/�?�?�<X|fҀ� �H�O :OJLOmOzI�J
! %@p1�O�O�O �O"3 __$_6_H_Z_l_ �n_�_�_�_�_@�_�_�_o"o\�e1o Vohozo�o�o�o�o�o �o�o
.@Rd`v���O5SK�0��8���?���F�4� X�H2OJ�AJ� [@G��A\O����(�O"�Oяb������p�O�z0  	� ��0p�Z�l�~�r_���9���ӟ���	��� $�C�7og� y���������ӯ��� 	��-�?�Q�c�u���𙿫����T1SV�GUNSPD%% �'%��2MO�DE_LIM �a9"ܴ2�	�� D-۵ASK_OPTION �9!�F�_DI EN�B  �5%f�B�C2_GRP 2�!�u#o2��XB��C����ԼBCCFGg #��*< #6���`�@I�4� Y��jߣߎ��߲��� ������E�0�i�T� ��x���������� ��/��S�>�w���+� t���u�����c��� 	B-f�.��4[  �������  02Dzh�� �����/
/@/ ./d/R/�/v/�/�/�/ �/�(���/?&?8?J? �/n?\?~?�?�?�?�? �?�?O�?4O"OXOFO hOjO|O�O�O�O�O�O �O__._T_B_x_f_ �_�_�_�_�_�_�_o o>o�/Voho�o�o�o (o�o�o�o�o(: Lp^���� ���� �6�$�Z� H�~�l�������؏Ə ��� ��0�2�D�z� h���To��ȟ���
� ��.��>�d�R����� ��z�Я������� (�*�<�r�`������� ��޿̿���8�&� \�Jπ�nϐϒϤ��� ���ϴ��(�F�X�j� �ώ�|ߞ��߲����� ���0��T�B�x�f� ������������� �>�,�N�t�b����� ������������: (^�v���� H���$HZ l:�~���� ���2/ /V/D/z/ h/�/�/�/�/�/�/�/ ?
?@?.?P?R?d?�? �?�?t�?�?OO*O �?NO<O^O�OrO�O�O �O�O�O�O__8_&_ H_J_\_�_�_�_�_�_ �_�_�_o4o"oXoFo |ojo�o�o�o�o�o�o �o�?6Hfx� �������v�&��$TBCSG_GRP 2$�u��  ��&� 
 ?�  Q�c�M���q��� �����ˏ��*�1��&8�d, ��F�?&�	 HCA;����b��?CS�B�I���<��V�>��ͪ�n��Ќ�ԝB��33Y3��Blt�������AÐ�fff�:��.�C����l�?����G�w�R���A&��̧�����@��I��-���
� X�u�@�R�����̻������	V3.0}0I�	mt7����*� �%��ֶY���@ff&� &�H�� N� �O�w  ����� �X�Ϙ�*�J21�'8���Ϥ�CFG -)�uB� E���+���d���#��#�I�W��pW� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ��������I�cp "4��gRw�� ����	-? �cN�r��&� �����/</*/ `/N/�/r/�/�/�/�/ �/?�/&??J?8?Z? \?n?�?�?�?�?�?�? O�? OFO4OjOXO�O �O`�O�OtO�O_�O 0__T_B_x_f_�_�_ �_�_�_�_�_�_,oo Poboto�o@o�o�o�o �o�o�o�o(L: p^������ �� �6�$�F�H�Z� ��~�����؏Ə��� �2��OJ�\�n���� ����������
� @�R�d�v�4������� ��ί����ү(�N� <�r�`���������ʿ ̿޿��8�&�\�J� ��nϐ϶Ϥ������� ��"��2�4�F�|�j� �ߎ����߀��� �� ��B�0�f�T��x�� �����������>� ,�b�P���������v� ������:(^ L�p�����  �$H6lZ |������/ �/ /2/h/�߀/�/ �/N/�/�/�/
?�/.? ?R?@?v?�?�?�?j? �?�?�?�?O*O<ONO OO�OrO�O�O�O�O �O�O _&__J_8_n_ \_�_�_�_�_�_�_�_ o�_4o"oXoFoho�o |o�o�o�o�o�o�/ $6�/�oxf�� ������,�>� ��t�b�������Ώ ��򏬏��&�(�:� p�^���������ܟʟ �� �6�$�Z�H�~� l�������دƯ���  ��D�2�T�z�h��� Jȿڿ������
� @�.�d�Rψ�vϬϾ� ���Ϡ������*� `�r߄ߖ�Pߺߨ��� �������&�\�J� ��n���������� ��"��F�4�j�X�z� |������������� 0B�Zl~(� ������, Pbt�D���8���   #� &0/"�$�TBJOP_GR�P 2*���  ?��&	H"O#,V,����� �z� =k%  Ȫ �� �� �$ �@ g"	 �C�A��&��SC���_%g!�"G���"k��/�+=��CS�?���?�&0%0CR  B4�'??J7��/�/?333�2Yx&0}?�:;��v 2R�1�0-1*20�6?��?20��7C�  �D�!�,� BL���OK:�Z�B_l  @pB@�� /s33C�1 �?gOO  A�zG�2jG��&)A)E�O�J;�}�|A?�ff@U@�1C�Z0zjO�Oz@ǰ��U�O�$ff�f0R)_;^;xCsQ?ٶ4)@�O�_tF��X_J\EU�_�V:�t-�Q(B�*@�Oo h�&-h$oZGLo6oDo ro�o~o8o�o�o�o�o 3�oRlVd(��V4�&`�q�%	V3.00m#Omt7A@�s*��l$!�'� E���qE���E��]\E�HF�P=F�{F�*HfF@D�F�W�3Fp?F��MF���F��MF��F��şF��F��=F���G�G.8��CW�RD3l)�D��E"���Ex�
E���E�,)FdR�FBFHFn� �F��F��M�F�ɽF�,
�GlGg!�G)�G=���GS5�GiĈ�;��
;�o��|& : @Xz�&/��&"�?��0�&=;-ESTP?ARS  (a �E#HRw�ABLEw 1-V) @�#R�7� � �R��R�R�'#!R�	�R�
R�R���!�R�R�R���RDI��`!��ԟ���
�r�Oz����� ����̯ޮ��Sx�^# <�����ÿտ��� ��/�A�S�e�wω� �ϭϿ�������;-w� {�_"��6��1�C�U� ��%�7�I�[���ҿNUM  �U`!� $  ���m���_CFG �.���!@H IM?EBF_TT}���^#��G�VE10m�H�z]�G�R 1/��O 8�" 2�� �A�  ��� ��������� �2�D� V�h�z����������� ��/
e@Rh v������� *<N`r� �����'/// ]/8/J/`/n/�/�/�/H�/r���_��t�@~��t�MI_CHA�NS� ~� !3DB/GLVLS�~�s��$0ETHERADW ?��w0�"���/�/�?�?l�$0R�OUTq�!�!��4�?�<SNMA�SKl8~�}1255.2E�s0OBOTO�s�t�OOLOFS_�DI}��%V9OR�QCTRL 0���#��MT�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo&l��OIo8omoq�PE_�DETAIJ8�JP�GL_CONFI�G 6�ᄀ�/cell/$�CID$/grp1qo�o�o/���?Zl~��� C���� �2�� V�h�z�������?�Q� ���
��.�@�Ϗd� v���������M���� ��*�<�˟ݟr��� ������̯@�}a�� �&�8�J�\���^o��c��`���˿ݿ�� �Z�7�I�[�m�ϑ�  ϵ����������!� ��E�W�i�{ߍߟ�.� �����������A� S�e�w����<��� ������+���O�a� s�������8������� '9��]o� ���F��� #5�Yk}������`�Us�er View ��i}}1234567890�//�,/>/P/X$� �cx/���2�U�/�/�/@�/??s/�/�3�/ b?t?�?�?�?�??�?�.4Q?O(O:OLO^OpO�?�O�.5O�O�O��O __$_�OE_�.6 �O~_�_�_�_�_�_7_�_�.7m_2oDoVoho zo�o�_�o�.8!o�o �o
.@�oagr� lCamera��o�� ��� �ޢE�*� <�N��h�z��������I  �v�)�� $�6�H�Z�l������ ����؟���� �2�Y��vP9ɟ~����� ��Ưد���� �k� D�V�h�z�����E�W� I5����� �2�D� �h�zό�׿������ ����
߱�W�ދ��X� j�|ߎߠ߲�Y����� ��E��0�B�T�f�x� ߁ulY��������� 
����@�R�d���� ������������W� i y�.@Rdv�/� ����* <N��W��i��� �����/*/</ �`/r/�/�/�/�/as9F/�/??1?C? U?�f?�?�?D/�?�?@�?�?	OO-O�j	�u0�?hOzO�O�O�O�O i?�O�O
_�?._@_R_ d_v_�_/OAO�p�{,_ �_�_oo)o;o�O_o qo�o�_�o�o�o�o�o �_�u���oM_q ���No���: �%�7�I�[�m�NE a����ˏݏ��� �7�I�[�������� ��ǟٟ����ͻp�%� 7�I�[�m��&����� ǯ�����!�3�E� 쟒�9�ܯ������ǿ ٿ뿒��!�3�~�W� i�{ύϟϱ�X����� H����!�3�E�W��� {ߍߟ�����������x����  �� L�^�p������������ ��    "�*�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/܄/�  
��( � �@�( 	 �/�/�/�/�/? ? 6?$?F?H?Z?�?~?�?�?�?�*2� � l�O/OAO��eOwO�O �O�O�O��O�O�O_ TO1_C_U_g_y_�_�O �_�_�__�_	oo-o ?oQo�_uo�o�o�_�o �o�o�o^opoM _q�o����� �6�%�7�~[�m� ��������ُ��� D�!�3�E�W�i�{� ԏ��ß՟����� /�A�S���w������ ��ѯ�����`�=� O�a�����������Ϳ ߿&�8��'�9π�]� oρϓϥϷ������� ��F�#�5�G�Y�k�}� �ϡ߳��������� �1�C�ߜ�y��� ����������	��b� ?�Q�c���������� ����(�)p�M�_q������0@� �������� ��#frh�:\tpgl\r�obots\m1�0ia4_7l.xml�Xj|��������.��/1/C/U/g/y/�/ �/�/�/�/�/�//? -???Q?c?u?�?�?�? �?�?�?�?
?O)O;O MO_OqO�O�O�O�O�O �O�OO _%_7_I_[_ m__�_�_�_�_�_�_ _�_!o3oEoWoio{o �o�o�o�o�o�o�_�o /ASew�� �����o��+� =�O�a�s����������͏ߏ�I ��<<  ?��4��,� N�|�b�������ʟ� Ο���0��8�f�L��~���������������(�$TPGL�_OUTPUT s9����� $�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ�@�ϳ�����$�����2345678901��� �2�D�V� ^����υߗߩ߻��� ��w����'�9�K�]���}g�������� o����1�C�U�g� ��u�����������}� ��-?Qc�� ������� );M_q	� ������%/7/ I/[/m///�/�/�/ �/�/�/�/?3?E?W? i?{??%?�?�?�?�? �?O�?OAOSOeOwO �O!O�O�O�O�O�O_��O� $$ Ӣ��OW=_o_a_�_�_ �_�_�_�_�_�_#oo Go9oko]o�o�o�o�o �o�o�o�oC5g}���������}@��"��? ( 	 iW� E�{�i�����Ï��ӏ Տ���A�/�e�S� ��w��������џ� ��+��;�=�O���s�����Ƹ  <<\ޯ�)�ͯ� )��M�_���ʯ���� <���ؿ��Ŀ� �~� $�V��BόϞ�x��� ��2ϼ�
ߤ���@�R� ,�v߈���p߾���j� ������<�߬�r� ���������� `�&�8���$�n�H�Z� �������������" 4Xj��R�� L����| Tf ��v�� 0B//�&/P/*/ </�/�/��/�/h/�/ ??�/:?L?�/4?�? ?n?�?�?�?�? O^? �?6OHO�?lO~OXO�O �OO$O�O�O�O_2_ __h_z_�O�_�_J_��_�_�_�_o.o��)�WGL1.XM�L�cm�$TPOFF_LIM Š|�p���qf�N_SVy`  ��t�jP_MON7 :���d�p��p2miSTRT?CHK ;���f�~tbVTCOM�PAT�h*q�fVW�VAR <�m\Mx�d  e��p�bua_DE�FPROG %��i%MAIN� P_p_REC�EPTOR|tb_DISPLAY�`��n�rINST_M�SK  �| >�zINUSE�p"ΕrLCK)��{QU?ICKMENM��toSCREl���~+rtpsc�t�)������b��_��S�Tz�iRACE_�CFG =�i�Mt�`	nt
?�~�HNL 2>�z���T{ zr@�R�d��v���������К�I�TEM 2?,�� �%$1234?567890�%�  =<�C�U�]��  !c�k�wp '���ns�ѯ5���� k������j�ů��� ����A�1�C�U�o�y� 󿝿I�oρ�忥�	� �-ϧ�Q���#�5ߙ� A߽�����e߳���� ��M���q߃�L��g� �ߋ����%�w� � [���+�Q�c���o� �������3��� {�;������G_�� ��/�Se.� I�m�� �=�a/3/�� ����k//�/�/ �/]/?�/�/�/?�/ u?�?�??�?5?G?Y? �?+O�?OOaO�?mO�? �?�OO�OCO__yO +_�O�Ox_�O�_�O�_ �_�_?_�_c_u_�_o �_Wo}o�o�_�oo)o ;o�o�oqo1C�oO �o�o��%��@[��Z��S��@��_��  �ے_� ����y
� Ï�Џ����UD1:\����q�R_GRP 1�A �� 	 @�pe�w�a���������ߟ͞�����ّ�>�)�b�M�?�  }���y�����ӯ ������	��Q�?� u�c���������Ϳ��	-���o�SC�B 2B{�  h�e�wωϛϭϿ��������e�UTORIAL C{��@��j�V_CONFIG D{����������O�OUTPUT� E{�����������%�7�I� [�m�������� ������%�7�I�[� m�������������� ��!3EWi{ �������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/��/??'?9?K? ]?o?�?�?�?�?�?�/ �?�?O#O5OGOYOkO }O�O�O�O�O�O�?�O __1_C_U_g_y_�_ �_�_�_�_�O�_	oo -o?oQocouo�o�o�o �o�o�_�o); M_q����� �yߋ����-�?�Q� c�u���������Ϗ� ��o�)�;�M�_�q� ��������˟ݟ� � �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i�{������� ÿտ���
��/�A� S�e�wωϛϭϿ��� ������+�=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� �����������1 CUgy���� ���	-?Q cu��������/�x��� $/6/ !/a/��/�/ �/�/�/�/�/??'? 9?K?]?�?�?�?�? �?�?�?�?O#O5OGO YOkO|?�O�O�O�O�O �O�O__1_C_U_g_ xO�_�_�_�_�_�_�_ 	oo-o?oQocot_�o �o�o�o�o�o�o );M_q�o�� ������%�7� I�[�m�~������Ǐ ُ����!�3�E�W� i�z�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'��9�K�]�o�~��$T�X_SCREEN� 1F8%  �}�~���������
����m&�� \�n߀ߒߤ߶�-�?� �����"�4�F��j� �ߎ���������_� ���0�B�T�f�x��� ���������� ��>��bt��� �3�W(: L^������ ��e/�6/H/Z/�l/~/�//�/�$U�ALRM_MSG� ?�����  �/���/�/)??M?@? q?d?v?�?�?�?�?�?��?O�%SEV  ��-EF�"EC�FG H����  ��@� � AuA   B���
 O���ŨO �O�O�O�O__&_8_�J_\_jWQAGRP �2I[K 0��	� �O�_� I_B�BL_NOTE �J[JT�G�l������g@~�RDEFPRO� �%�+ (%C�OLOCA_ME�SA_IRVISION�_%OVoAo zoeo�o�o�o�o�o�o��o@�[FKE�YDATA 1K<�ɞPp jG���_������z�,(����([ INST ]'�<)�v@NCELS�~���NDIRECT���� ES  S�TEP��*�[E�DCMDB���ORE<�FO��C� U�<�y�`�������ӟ ����	��-��Q�c�� ��/fr�h/gui/wh�itehome.pngd�����Ưد�ꯀ{�inst����/�A�S�e��� � FRH/FCG�TP/wzcancel�����˿ݿ��~� �direc��(�:�L�^�p���yes�ϭϿ����������{�edcmd��3�E�W�i�{����{�arwrg ϲ���������y�� )�;�M�_�q���� �����������%�7� I�[�m��������� ��������3EW i{����� ��/ASew ��r������ /!/(E/W/i/{/�/ �/./�/�/�/�/?? �//?S?e?w?�?�?�? <?�?�?�?OO+O�? OOaOsO�O�O�O8O�O �O�O__'_9_�O]_ o_�_�_�_�_F_�_�_ �_o#o5o�_Goko}o �o�o�o�oTo�o�o 1C�ogy�� ��P��	��-� ?�Q��u����������Ϗj�܋�u� ܏�(�s��Q�c�r��,I���A�POI�NT ER��9� ?OOK T ßğ�  NDIREC�T�� CHOI�CE]��TOUCHUPG�H�s� ��~�����߯�د� ��9�K�2�o�V�����茿ɿ��whi?tehome���� �2�D�V�	�poin�ߍϟϱ�����`��look��#��5�G�Y���i/indirec|Ϙߪ���������choic���� �2�D�V�h��k��touchup�ߠ���������g��arwrg ��"�4�F�X�j�a��� ����������w� 0BTfx�� �����,> Pbt���� ��/�(/:/L/^/ p/�//�/�/�/�/�/  ?׿�/6?H?Z?l?~? �?�/�?�?�?�?�?O �?2ODOVOhOzO�O�O -O�O�O�O�O
__�O @_R_d_v_�_�_)_�_ �_�_�_oo*o�_No `oro�o�o�o7o�o�o �o&�oJ\n ����E��� �"�4��X�j�|��� ����A�֏����� 0�B�яf�x������� ��O������,�>��ټL������u�����q���ͯ��,������"�	� F�X�?�|�c������� ֿ������0��T� f�Mϊ�qϮϕ����� �����,�>�?b�t� �ߘߪ߼�˟����� �(�:�L���p��� �����Y��� ��$� 6�H���l�~������� ����g��� 2D V��z����� c�
.@Rd �������q //*/</N/`/��/ �/�/�/�/�/�//? &?8?J?\?n?�/�?�? �?�?�?�?{?O"O4O FOXOjO|OSߠO�O�O �O�O�OO_0_B_T_ f_x_�__�_�_�_�_ �_o�_,o>oPoboto �oo�o�o�o�o�o �o:L^p�� #���� ��� 6�H�Z�l�~�����1� Ə؏���� ���D� V�h�z�����-�ԟ ���
��.���R�d� v�������;�Я��� ��*���N�`�r���Ж������@���>�@������ 	��+�=��,)�n� !ߒ�y϶��ϯ����� �"�	�F�-�j�|�c� �߇����߽������ �B�T�;�x�_��� �O��������,�;� P�b�t���������K� ����(:��^ p����G��  $6H�l~ ����U��/  /2/D/�h/z/�/�/ �/�/�/c/�/
??.? @?R?�/v?�?�?�?�? �?_?�?OO*O<ONO `O�?�O�O�O�O�O�O mO__&_8_J_\_�O �_�_�_�_�_�_�_�� o"o4oFoXojoq_�o �o�o�o�o�o�o�o 0BTfx�� ������,�>� P�b�t��������Ώ ������(�:�L�^� p��������ʟܟ�  ����6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z����� -�¿Կ���
�ϫ� @�R�d�vψϚ�)Ͼπ��������*�`�,��`���U�g�y�Qߛ߭߇�,���ߑ����&�8� �\�C���y��� ���������4�F�-� j�Q���u��������� ���_BTfx �������� ,�Pbt�� �9���//(/ �L/^/p/�/�/�/�/ G/�/�/ ??$?6?�/ Z?l?~?�?�?�?C?�? �?�?O O2ODO�?hO zO�O�O�O�OQO�O�O 
__._@_�Od_v_�_ �_�_�_�___�_oo *o<oNo�_ro�o�o�o �o�o[o�o&8 J\3����� ��o��"�4�F�X� j��������ď֏� w���0�B�T�f��� ��������ҟ����� �,�>�P�b�t���� ����ί�򯁯�(� :�L�^�p�������� ʿܿ� Ϗ�$�6�H� Z�l�~�Ϣϴ����� ����ߝ�2�D�V�h� zߌ�߰��������� 
��.�@�R�d�v�ﴚ�qp���qp���������������,	N�r� Y������������� ��&J\C�g �������" 4X?|�m� ����/�0/B/ T/f/x/�/�/+/�/�/ �/�/??�/>?P?b? t?�?�?'?�?�?�?�? OO(O�?LO^OpO�O �O�O5O�O�O�O __ $_�OH_Z_l_~_�_�_ �_C_�_�_�_o o2o �_Vohozo�o�o�o?o �o�o�o
.@�o dv����M� ���*�<��`�r� ��������̏���� �&�8�J�Q�n����� ����ȟڟi����"� 4�F�X��|������� į֯e�����0�B� T�f�����������ҿ �s���,�>�P�b� �ϘϪϼ������� ���(�:�L�^�p��� �ߦ߸�������}�� $�6�H�Z�l�~��� ����������� �2� D�V�h�z�	��������������
�}�����5@GY1{�g,y �q���< #`rY�}�� ���/&//J/1/ n/U/�/�/�/�/�/�/ �/ݏ"?4?F?X?j?|? ���?�?�?�?�?�?O �?0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�_�_'_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o $�oHZl ~��1���� � ��D�V�h�z��� ����?�ԏ���
�� .���R�d�v������� ;�П�����*�<� ?`�r����������� ޯ���&�8�J�ٯ n���������ȿW�� ���"�4�F�տj�|� �Ϡϲ�����e���� �0�B�T���xߊߜ� ������a�����,� >�P�b��߆���� ����o���(�:�L� ^�������������� ��}�$6HZl ��������y  2DVhzQ��|�Q�����������,�/./�/R/9/v/ �/o/�/�/�/�/�/? �/*?<?#?`?G?�?�? }?�?�?�?�?OO�? 8OO\OnOM��O�O�O �O�O�O�_"_4_F_ X_j_|__�_�_�_�_ �_�_�_o0oBoTofo xoo�o�o�o�o�o�o �o,>Pbt� ������� (�:�L�^�p�����#� ��ʏ܏� ����6� H�Z�l�~������Ɵ ؟���� ���D�V� h�z�����-�¯ԯ� ��
����@�R�d�v� �������Oп���� �*�1�N�`�rτϖ� �Ϻ�I�������&� 8���\�n߀ߒߤ߶� E��������"�4�F� ��j�|������S� ������0�B���f� x�����������a��� ,>P��t� ����]� (:L^���� ���k //$/6/ H/Z/�~/�/�/�/�/h�/�/���+������?'?9=?[?m?G6,YO�?QO �?�?�?�?�?OO@O RO9OvO]O�O�O�O�O �O�O_�O*__N_5_ r_�_k_�_�_�_�_�� oo&o8oJo\ok/�o �o�o�o�o�o�o{o "4FXj�o�� ����w��0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� ����(�:�L�^�p� �������ʯܯ� � ��$�6�H�Z�l�~��� ���ƿؿ���ϝ� 2�D�V�h�zό�ϰ� ��������
���_@� R�d�v߈ߚߡϾ��� ������*��N�`� r����7������� ��&���J�\�n��� ������E������� "4��Xj|�� �A���0 B�fx���� O��//,/>/� b/t/�/�/�/�/�/]/ �/??(?:?L?�/p? �?�?�?�?�?Y?�? O�O$O6OHOZO�$U�I_INUSER  ���{A��  �[O_O_MENH�IST 1L{E�  (� �@��(/S�OFTPART/�GENLINK?�current=�menupage?,148,2�O_�_1_C_�O�O,19�1,1 ARRA�_ESTEIRA@~P�_�_�_�_�0)X_�j_63}QLACE0�_o.o@oK_�_�J54o�o�o�o�o�0	'`orn7}Q/�AS�_�gedit�BMAIN	����� �9hz~C�OLOCA�@SA�_IRVISIO��3�E�W��o�o�B2�3#�����ʏ܏�0���0�A����"�4�F�X�j� �������� şן�x���1�C� U�g�����������ӯ ������-�?�Q�c� u��������Ͽ�� ���)�;�M�_�qσ� ϧϹ��������� %�7�I�[�m�ߑߔ� ������������3� E�W�i�{������ ����������A�S� e�w�����*������� ����=Oas ���8��� '�0]o�� ������/#/ 5/�Y/k/}/�/�/�/ B/�/�/�/??1?C? �/g?y?�?�?�?�?P? �?�?	OO-O?O�?PO uO�O�O�O�O�O^O�O __)_;_M_8�O�_ �_�_�_�_�_�Ooo %o7oIo[o�_o�o�o �o�o�o�ozo!3 EWi�o���� ��v��/�A�S� e�w��������я� �����+�=�O�a�s��^[�$UI_PA�NEDATA 1�N������  	�}�c/frh/cg�tp/flexd�ev.stm?_�width=0&�_height=�10ԐŐice=�TP&_line�s=3Ԑcolu�mns=4Ԑfo�nܐ4&_pag�e=doubŐ1���\V)prim#�L�  }O�s���0������ͯ )ϯ� گ���;�M�4�q�X� ������˿������%�\V�� �E�  �N�"]�d��ɟ۞2�����2/�-�dual ����_��"�4�F�X� j�ώ�u߲��߫��� �����B�)�f�M�`������3� G�O8�����*�<� N�`�����Ϩ����� ����i�&8\ C��y���� ��4Xj=� ���������� �� /S$/��H/Z/ l/~/�/�/	/�/�/�/ �/�/ ?2??V?=?z? a?�?�?�?�?�?�?
O }�@OROdOvO�O�O �?�O1/�O�O__*_ <_N_�Or_Y_�_}_�_ �_�_�_�_o&ooJo 1ono�ogo�oO)O�o �o�o"4�oXj �O������O ��0�B�)�f�M��� �����������ݏ� �>��o�o������� ��Ο��3��w(�:� L�^�p���韦����� ܯï ����6��Z� A�~���w�����ؿ� ]�o� �2�D�V�h�z� Ϳ�����������
� �.ߕ�R�9�v�]ߚ� �ߓ��߷������*��N�`�G����	��������������"�) ��G���6�s������� ����4������� K2oV���� ����#������$UI_POSTYPE  ��� 	 �/�UQUICKMEN  d�s�WREST�ORE 1O��  �	�� /#���m+/T/f/x/�/�/?/ �/�/�/�/?�/,?>? P?b?t?/�?�?�?? �?�?OO(O�?LO^O pO�O�O�OIO�O�O�O  __�?_1_C_�O~_ �_�_�_�_i_�_�_o  o2o�_Vohozo�o�o I_So�o�oAo�o. @Rd���� �s���*�<��o I�[�m������̏ޏ �����&�8�J�\�n���������ȟڟ�S�CRE�?��u1sc��u2�3�4�5*�6�7�8��wTAT`� �<�MUSER������ks���3��4���5��6��7��8���UNDO_CFG Pd����U�PDX�����None���_INFO 1Q�5<��0%��W� ��E���i�������� �տ���:�L�/�p����eϦύ)�OFF?SET Td@���{������	�� -�Z�Q�cߐ߇ߙ��� �������� ��)�V� M�_�q�۹������
���t��)�WO_RK U4������A�S��ψ�UFR?AME  ����&�RTOL_AB�RT��$���ENB�����GRP 1V���Cz  A���+=O@as�����U�������MSK  h�<���N��%4���%��)��_EV�N�����>�2�W��
 h���UEV��!td�:\event_�user\-�C�7���}�F��S�P��spot�weld�!CA6����! �Z/�/:'�H/~/l/ �/�/�/�/-?�/Q?�/ ? ?�?D?�?h?z?�? O�?)O�?�?OqO`O �O@ORO�OvO�O_�O��O7_�O[__Z]Wf+�2X����8V_�_�_ �_�_o�_,o >oobotoOo�o�o�o �o�o�o�o:L�'p�]�����$VARS_CO�NFI�Y�� F�P{���|CCRG�\��>�{�ut�D� BH� Ypk�a�C�� ���}�?���C,&Q=���ͩ�A �MRv2b���	�}�	��@�%1:� SC130EFG2 *����{����Y�X� �5}������A@k�C�F� w�Q�[���|�@���������T��ā�\�ϟ �\� B���;�e�@� ǟ`�����S�����̯ ���ۯ�&�}��\��G�Y���E���ȿ�TCC�c
���������pGF�pgd���-�23456789017�0?��ׁ$���4�v�@Nm�� ��϶�BW������i�}�:�o=LA�څ�6�@�6� ͿZ���i�7����(��W���-�]�X�jĈ� �ߕϳϹ�������� �%�7�I�r�m�ߨ� �ߵ����������8� 3�E�W������}��� ����������/�A��S�e�w��MODE���t �RSL�T e�|k�%" zς��;�1��d���`��SELE�C��c��	IA�_WO�Pf �� W,	�	������G�P� �����RTS�YNCSE� ���$�	#WINURLg ?*ـ�;�\/n/�/�/�/�/�uI�SIONTMOU8���A# ��%��gSۣ�Sۥ�P�� FR:�\�#\DATA\��/ �� M�C6LOG?  � UD16EX�@?\�' B@� ���2T1G�abriel_Fariak?P5�?�?������ n6  ���GV�2\�� -��5�� �  ��Z�@U0>58TRAINj?��4*B{Rd_Cp��D #`{2��'$t�"��h#� (� kI�Mw��O�O�O�O�O 1__U_C_]_g_y_�_��_�_�(STA� i���@��o0oI:$�obo�%_GE�jv#��~@ �
��\��btgHOMIN��kSۮ��`�P2,,��CWǖB�veJMPERR {2l#�
  Qo I:��"�4Fwj |����������&%S_g0REr�m�^۴LEXd�n�1-ehoV�MPHASE  ��e׃BޱOF�F _ENB  ��$VP2�$o/Sۯ��x�c C;�@ �@�;����?s33'D*AA ��]� ��0ޱ�`r}�XC��܅���p\A-۟E �� ����#�5������� ������}�������� ��c�X���A����� ϯ�+��߿��M� B�q���xϊϹ���� ��������7�I�;�m� b�)ߣ�Eߓߡ߳��� ��3���W�L�{ߍ� �ߑ���������� /�$�6�e�W���c�y� ������������� O���?M_q��� ����'9�= 7Is����� �/m/%/3/E/�s�TD_FILTuE�`s�k �x2�`����/�/�/�/ �/	??-???Q?�6�/ ~?�?�?�?�?�?�?�?�O OoiSHIFTMENU 1t}<5�%5�~O)�\O �O�O�O�O�O�O�O'_ �O_6_o_F_X_�_|_��_�_�_	LIV�E/SNAP�S?vsfliv���_��z`ION �ҀU
`bmenu &o+o�_�o�oV"<E�uz��4IMO�v����zq�WAIT�DINEND  a�ec��b�fOKوNOUT�hSD�yTIMdu��o|G�}#�{C�z�b�z�xRELE���ڋxTM�{�d=��c_ACT`و���x_DATA �wz���%  E�GA_BARRA�_ESTEIRAx�o6Ex�RDIS
`~E��$XVR�a�x�n�$ZAB�C_GRP 1yvz��� ,��2̏.MZD��CSKCH�`z���aP@��h@�IP�b{'���şן�[��MPCF_G 1|'���0�r�8�d�� �}'��p�s�� 	(���  �<l0  ���X;?�  4
�D���5�X=�������4�
C�����?���C�8�D��w�>w�@2�����<�X���gs��`8��v>������ɯ ۯ�����o���w�ܴ�� /��3�������B� ˿ݸĸ+��	���1�?�i�����x�3ɟ]�6��y��W����3ɝ�+��C|3��7�i��0��?�׌����'>�
a�������Rw>C��:�[�	��`~�����_CYLIND�~!� Р? ,(  *.�?���+�h�Oߌ�s�  ��������(�	�x�-� �&�c�߇����� ��j�P����)��~�0_�q��� �2�'��� �&��������@��&��I��c�A���SPHER/E 2����� �����A�T/ A��e���� ��/N`=/� a/H/Z/�/��/�/�/6�ZZ� ��f