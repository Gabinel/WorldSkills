��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� � P�COUPLE,  o $�!PPV1OCES0�!H1�!��PR0�2	 � $SOFT��T_IDBTOT_AL_EQ� Q1�]@NO`BU SPI�_INDE]uEX�BSCREEN_��4BSIG�0�O%KW@PK_F�I0	$TH{KY�GPANEhD� � DUMMYE1d�D�!U4 Q�!RG1R�
 � $TIT1 d ��� 7Td7T� 7TTP7T55V65V75V85V95W05W>W�A�7URWQ7UfW1pW1
zW1�W1�W 6P!�SBN_CF�!-�0$!J� ; |
2�1_CMNT�$FLAGS]n�CHE"$Nb�_OPT�3�(C�ELLSETUP�  `�0HO��0 PRZ1%{cM�ACRO�bREP	R�hD0D+t@��bl{�eHM MN�yB
1�UTOB �U�0 �9DEVIC4ST	I�0�� P@13�r�`BQdf"VAL�#ISP_UNI��#p_DOv7IyFR_F�@K%D13�x;A�c�C_WA?t��a�zOFF_@N.�DEL�xLF0q8�A�qr?q�pF�C?�`�A�E�C#��s�ATB�t�d��MO� �sE �� [M�s��2�R;EV�BILF��1�XI� %�R � � OD}`j�_$NO`M� +��b�x�/�"u��� ����!X�@D�d p E R�D_Eb��$F�SSB�&W`KBD�_SE2uAG� G
�2 "_��B�� V�t:5`ׁQC �a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR�B�IGALLOW�� (KD2�2�@VAR5�d!�AB �e`BL[@S � !,KJqM�H`S�pZ@�M_O]z����CFd X�0G�R@��M�NF�LI���;@UIR�E�84�"� SWIYT=$/0_No`S�"�CFd0M� =�#PEED��!��%`���p3`J3tV�&$E�..p`L�>�ELBOF� ��m��m�p/0��CP�� F�B����1���r@1J1E_y_T>!Բ�`��g����G� �0WARNMxp�d�%`��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqM��� R�r$ORIأ.&ӧRT�SF\g CHGV0I�Ep�T��PA�I{��T�!��� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5��6�7�8�9��4��x@�2 @.� TRQ��$%f��4ր����_U����z��Oc <� �����Ȩ3�2��LL�ECM�-�MULTIV4�"$��A
2q�CHILD>�
1���z@T_1b  4� STY2�b4�=@�)24����@��� |9$��T��A�I`�E��eTOt���E��EXT����ᗑ�B��22(�0>��@��1b�.'��}!�A�K�  �"K�/%�a��R���N?s  =�O�!M���;A�֗�M�� 	��  =�I�" �L�0[�� R�pA��$JOBB�����ނ�TRIGI�# dӀ����R�-'r0��A�ҧ��_M��b7$ tӀFL6�BsNG�A��TBA�  ϑ�!��
/1�À�0���R0�P/p ����%�|��Bqh@W�
2JW�_RH��CZJZ�_zJ
?�D/5C�	�ӧ�t�@��Rd&�������ȯ�qGӨg@N�HANC��$LG /��a2qӐ� ـ@��!A�p� ���aR��0>$x��?#DB�?#3RA�c?#AZt@�(p.�����`FCT��ƕ�_F࠳`�SM��!I�+lA�%` � ` ���$/�/����[�a��M�0\��`l��أHK��AEs@�͐�!�"W��N� SbXYZW�`�"�����6	��I���'  . I�I��2�(p�STD�_C�t�1Q��US�TڒU�)#�0U�[�%?IO1��� _Up�q�* \��=�#AORzs8Bp�;�]��`O6  RSY�G�0�q^EUp��H`�G�� ��]�DBPX�WORK�+* $SKP_�p��A��TR�p , �=�`����Z m�O1D3��a _C"�;b�C� �GPL:c�a�tDőS�D�W�3B�b����P��P &)DB�!�-�B APR��
I�Ja3��. /�u������K�LuY/�_�����0�_���PC��1�_���~�EG�]� 2�_�SVP�RE.��R3H �$C��.$L�8c/$uSނz IkI3NE�WA_D1%�ROyp�������q0�c7 t@�fPA���?RETURN�b��MMR"U��I�C�Rg`EWM@�SIGNZ�A ��|�e� 0$P'��1$P� m�2�p�p'tm�+pD��@ �'�bdNa)r�GO_AW ��@4ؑB1I�CSd�(�KCYI�4���`1w��qu��t2�z2�vN��}��E}sDEV�Is` 5 P �$��RB��I�wPk��I_BYȧ��"�T7Q�tHN{DG�Q6 H4���1�w��$DSBLC��o��vg@��|tL��7O�f@]���3FB���FEra8��ׂ�t}s���8> pi�T1?���MCS����fD �ւ[2H� W ��EE���%F����t����9 T�p��x�NK_N:�����UZ��L�wHA�vZ' ~�2���P~r�q7w: �=MDLn��9�ጂٱh����! e����J��~� +����,�N�D����3���ՒG!aqSL�Ad�7;  ��INP��"�����}q_ V�4<�06`C� �NU��  D�L�ק��SH!�7=BM��q���ܢӢ����g���>P +$ٰ�٢��^��^�Y�FI B�\��Ă��'A	'AW�l�NTV��]�V\~�X�SKI�#T� ��a�ۺ�T1J�3:39_�P�SAFN����_SV�EXCSLU��N@�DV@�Ll @�Y����S�H�I_V
0\2PPL5YPRo�HIM�T��n�_MLX��pVORFY_�Cl�M��gIOC�UC_� �����O�q�LS(�0v�FT4Q���)��@P�E$�t��A��CNFt�6եup��pm�4ACHD��o������AFC C	PlV�TQTP?�� ί� ?`�@TA��@�0L@ ��N���]� @����T��T! S����te@{R�A DO�� w23���!n��	_1�#�H!�̔�΀�K��B�2��MAR�GI�$���A ���_SGNE�C;
$�`�a^aR0 ��3��@ B��B��ANNUN�P?����uCN@�`%0��`��� ���BEFc@]I�RD @Q�F���4OT�`�sFTӠHR,Q��CQ0�M��N�I|RE�����A�W���DAY=CLOCAD�t;T|�<S5}�EFF_AXI��%F`1QO3O��Eq���@_RTRQ�E�G����0RQ
�2Evp ��|��F�0f�R0 �tM��AMP�E<� H 0�`œ^��`Ds�DU�`��v�BCAr� I?��`N ErIDLE_PWRI\V!n0�V�wV_[ |�� ��DIAG�5J�o 1$V�`SE�3TQl�e��P�l�^E_��Y�VE6� �0SWH�q (� �b|�Gn�3OHxPPHZ�IRAl�B�@�[� �a�b�1�w3�O  � ��v�|�I�0 ��pRQDW�MS-�%AX{6Y�LIFE�@�&�MQy�NH!Q%��F#�C����CB0�mpNr$�Y @�aFLAl�f��OV0]&HE��>l�SUPPO�@u��y��@_�$��!_�X83�$gq�'Z�*W��*B1�'T�#`�k2XYZáY�Y2D8CY`T@�`N�����f� �C�I2��IC�TA�K `�pCACH�ӫ�3�����I��bNӰUFFI� \��@��;T��r<S6CQ.�MSW�5�L 8	�KEYI7MAG�cTMLa���*Ax�&E���B��OC�VIER-aM ���BGL����y�?G� 	��П4N�m:�ST�!�B P�D,P�D��D��@�EMAI䐔a��M��r�FAUL|RO bB�c�� spUʰMA�"`T'`E�P< �$S�S[ � ITw�BUF�7y��7r�tN[�LSUB1T��Cx�o�R�tRSAV|U>R'c2�\�WT���P�T�*`S�n�_1PbU���YOT(�bK��P��M��d����WAX��2��XX1P��S_GH#
���YN_���Q <�Q�D��0���M��� T�F�`�|�\�DI��EDT�_Pɰ:�R��b�G�RQM�&��Jq�a����׀��Fs� S (�SVqpB��4��_�.��a��T�� �@���B�SC_R]1IK>B'r��$t�R"A#u�H�aDS�P:FrP�lyIM@|Sas�qz��a� U>wh� <1%sM�@IP��0s��0`tTHb0ЃdTr��T`asHS�c�CsBSCʴq0� V`�����S�_D��/CONVE�G���Hb0^v1PFHy�dCs�`&a?ASC���s�MERg��aFBC�MPg��`ET[� �UBFU� DU�%P�D�:12�CD�Wy�p�P�CG�[@N	O6�:�V� ��� �R��P���C������w��A��`��W/H *�LƠ�C c�W����Y�賂��� ��q�|���A*��7}�8}�9}�H T���1��1��1��U1��1ʚ1ך1䚕1�2��2����2���2��2��2ʚ2�ך2�2�3��3R��3����3��3��U3ʚ3ך3�3�94��QEXT[�X[b�H``t&``z�k`t˷$���FDR�/YTPV��RpK"	��K"REM*9F��]"OVM:s/ŽA8�TROV8�D�T�PX�MXg�INp8ɉ W��INDv�BH2
�ȕ`K ^`G1a �a��@Q%7Da��RIV��u"]"GE[AR:qIO.K(�H4N�`���,(�F@|� I3Z_MCM<0.K! �F� UT����Z ,�TQ?� b�y@t�G?t�E |�.�>Q�����[ �Pa�� RI�E��UP?2_ \ �@=S#TD	p<TT����p�����a>RBACUbG] T��>R�d)�j�%C�E��0��IFI���0��i�{�4�PT�T��FLUI�D�^ �?0gHPUR �gQ�"�r�a�4P�+ I�$��Sd�k?x��J�`CO�P��SVRT��N�x$�SHO* ��CAS�S��Qw%�pٴBG_%��3���<�FORC�B��^o�DATA��_�BKFU_�1�bb�2�a�m=mm�b0��` �|��NAV	`)������$�S�Bu#?$VISI���2SC	dSE������V��O�$&�B�K�� ��$PO���I��FM�R2��a  ��	��`#��@&�8�O� (�_��9��+IT_^�ۄ�)M�����DGC{LF�DGDY�LD����5Y&��Q$RY�M됇CbN@{	? T�FS�P�D�c P��W�cK �$EX_WnW1P%`]��"X3�5�s�G+�d ���ָ�SWeUO�DE�BUG��-�GRt��;@U�BKU���O1R� _ P�O_ )�����M���LOOc>!SM E�R�a��u _E� e >@�G_�TERM`%fi'��ORI�ae gi%y�SM_�`>Re !hi%V�(ii%3�UP\Bj� -����e��w#� f���G�*ELTOr�A�bF�FIG�2��a_���@�$�$g$wUFR�b$�01R0օ� OT_7F��TA�p q3NST��`PAT�q�0�2P'THJ�ԀE�@�c3ART�P'58�Q�B�aREL�:�aSHFT�r�a�1�8E_��R��у�& � 	$�'@i�
����sN@bSHI�0�Uy�= �QAYLO�p� Oaq�����1����pERV��XA��H�� m7�`�2%�P�E3�P��RC���ASYM�a��aWJ07����AE�ӷ1�I��ׁUT@�`Oa�5�F�5P�sXu@J�7FOR�`M # �O!k]��`5&�0L0��`HOL ;l �s2T�����OC1!E��$OP��qn����$�����$��PR�^��aOU��3e���R�5e�X�1 �eo$PWR��IMe�BR_�S�4�� �3��aUD��k�Q�dm���$H�e!�`AWDDR˶HR!G�20�a�a�apRR��[�n H��S����%���e3��e���e��SE���z�HS�MNu�o���Pªq��0OL�s߰`ڵ<�I ACRO��&1��ND_C�s��A<fdK�ROUP��R!_�В� �Q1|�= �s���y%��y-��x�� �y���y>�=A�����AVED�w-��uy&sp $�І�P_D�� ��'rP�RM_���!HT�TP_�H[�q (ÀOBJ��b �[$˶LE~3��>\�r � ����J��_��TE#ԂS�P�IC��KRLPiHI�TCOU�!��L ���PԂ������PR���PSSB�{�JQUERY_FLAvs��@_WEBSOC����HW�#1��s��`<PINCPU(���O���g������d��t��O� �IwOLN�t 8��yR��$SL!�$INPUT_�U!$`��P �G֐SL.���u���2�.��C��B��IOa�F_AS:=v�$L+ਇ+�A��bb41�����Z@HYʷ�����#qe�UOP:w `v�ϡ˶�¡�������"`PIC`����� �	�H�IP_ME���v�x Xv�IP�`(�R�_N�p�d����Rʳp�ױQrSaP �z�C��BG(��� ��M�Av�y lLv@CTApB��AL TI�3UfP_ ۵�0�PSڶBU_ ID � 
�L � `�Q0��L��0z)�����ϴ�NN�_ O��I�RCA_CNf� �{ �Ɖ-�CYpEA������� �IC�ǫ�tpR�=Q�DAY_
��NTVA�����!��5�����SCAj@��CL��
����
���v�|`5�VĬ2b�l�N_�PACV�n�
���w�})� T��S�����
��e����T� 2| Ր�� �v�~��֣�ذLAB1��_ �חUNIX��ӑ ITY裪��e~�p�� ���<)���R_U�RL���$A;qEAN ���s`vsTeqwT_U��m�J��X�M�$���E��"��R祪�� A�,�2��JH���FLy���= 
���
�UJ]R|U� ���F��6G��K7��D>�$�J7�s��J8*�7����3�E�7��&�8�\�)�APHI�Q4�y�DkJ7Jy8R��L_KE'�  �K͐L}MX� � <U��XRi�����WATCH_VAZqu@Aស�FIEL`��cy�n���:� � u1VbwPCTX�j��Y �LGE���� !��LG_SIZ΄�[8Zm�ZFDeIYp1! gXb ZW �S`� 8�m��� �b ���A�0_i0_CM c3#�*'FQ1�KW d(V(Bbpo pm�p� |Io�1 pb p�W RS��0  M(C�LN�R�۠-�DE6E3��� �c�i���PL#�7DAU"%EAq�͐�T8". GH�R��y��BOO�a��3 C��F�ITV�l$�A0��RE���(SCRX����D&�ǒ�qMARGI�Sp�,@����T�"�y�S���x�W�$y�$��JG=M7MNCHt�y�FN��6K@7r�>9�UFL87@L8FWDvL8HL�9STPL:�VL8"�L8s L8RS"�9HOPh;��C9D�3 R��}P�'IUh�`4@�'�5$ ��S2G09�pPOWG�:�%�3,�64��N9EX��TUI>5I� �ӌ���� �C3�C<0'�,�o�:��&�@�!NaqvcAcNAy��Q�AI]�8gt7Ӝ�DCS���c�RS�cRROXXOdWS��ÂRoXS{X�(IGNp 
Ђ=10 ��[T�DEV�7LL���CZ!*�C �	 8�Tr$f/蛒����Z�3A�a�	 W�h萦�Oqs�S1Je2Je3Ja��BSPC G� �ƋG`-T� �%��Q�T�r@�&E�V�fST�R9 YBr~�a �$E�fC�k�g��f	v��CB� L����� �� u�xs뀔�g�q�jt:��!�#_ ����ʐv�#Ӡ �s �M�C�� ���C�LDP᠜�TRQ�LI ���y�tFL ���rQ��s5�D���w�~�LD�u�t�uOR�G���1�RESERV��M���M�Œ�C�s��� � a	�u�5�t�uSV���p��	1�����RCLMC��M�_�ωxА��: MDBGh��I����$DEBUGMAS������JU�$T8P��EF��d�
�MFRQ~Ҥ� � K	�HRS_RU��bq��A��$EFRE�QUu!$0YOVER�k��f��PU1EFI�%�Gq�� �6�Y�z��� \����E�$U��`��?��
�P)SI`��	��CA ���ʲ�σUY�%�?�( 	��MISC��� d��aRQ���	��TB� � 1���A��AX���|����EXCESg��d�M�H�9��u���9d�SC�` O� H�х�_��@���������pKE�a��+�� &�B_, �FLICBtB� QoUIRE CMOt�QO���r�LdpMD�� �p{!��5b����ND!��I�!���L �D;
$�INAUT�!
$R#SM�ȧPN����C�PSTLHᗻ 4U�LOC�fR�I"��eEX��ANqG.R.���ODA]���q��� �RMF0����icr�@mu8���$�SUPiu��FX��IGG! � ���cs�F� cs
Fct��ޒ�b5��` E��`T�5�tC��g�#TI��7�M���7� t��MD���A)��XP��ԁ��H��.���DIAa��Ӻ�AW�!��0af���D@#�)֡O�㥀��� -�CUp V	����.����!_��� ��{`�c������� |�P|��0� ��P�{�KEB��e-$qB��o�=pND2ւ�����2_TXltXGTRAXS������LO: ����}� ���C�.�&���RR2h���� -�!A�� ?d$CALI����GFQj�2F`RIN�bn�<$Rx�SWq0ۄ���ABC�ȇD_J��{�q��_�J3��
��1SPH, �q�P����3��(H�9pq�#J�34n���O�QIM�M�CSKP�zb7?SbJ+�M�Qb�y8����_AZ��/��EL�Q.ցOC�MP��N�� RTE�� �1�0 ����1��@ ZScMG�0����JG�p�SCLʠ��SPH�_�PM��f��q��u�RTER��n��Pk�_EP�q�`A0� �cM��DI�Q�23UdDF  쀐�LW�VEL��qINxr�@�_BALXP.��Y/�J�0�'$Q�IN���B]�C�9%�".�8!:6p_T� �F%a"�6#a!��k)�Q�DHʠ��\�9`�$Vw��_�A$�=����&A$���S�h��H ��$BEL� m��_oACCE� 	8<�0IRC_�q��@�NT��c$SPSʠ�rL��� M4�s9 .7��GP/6��9�7$3�73S2T�͡_Ga�"�0�1��8�17_MG}�DD�1���FW�p��3�5$3�2�8DEKPPA�BN[7ROgEE �2KaBO�p�Ka���1�$USE_tv�SP��CTRT�Y4@� �� <qYN�g�A�@�FR �ѢAM:�N�=R�0O�v1�DINC(��B�4����GY��ENC�L���.�K12��H0IN¿bIS28U��ONT|�%NT23_���fSLO���|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1��M�PERCH  �S��� �W���SlщR ��l����E�0�0P	AS2EeL�DP7�O�NUЉZ�f�VTRK�RqAY"�?c��a S2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gBT��DUX �2S_BC?KLSH_CS2Fu :��V���C-�esRoz|�A�CLALMJTp@��`� �uCHKe |����GLRTYp� ��8T��5���_�ùT'_UM3��vC3��1�Z���LMT��_ALG��%���0�E*� K�=�)�@5F�@8 9��Nb��)hPC�Q)hHpТ��5�uCMC��\�0�7CN_��N��L�;SF�!iV�B���.W���S2/�ĈCAT�~SH�Å��4  V�q/q/V�T1�f�0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e��R� @B�_Wu�d@�!a��#`��#`�Ih�Iv�I�#F��S�:X��I�0VC00��֢1ܮ�0�⦇JRKܬ!��<�D�BXMt�<�M�_sDL�!_bGRVg�``��#`��#A�H_%�8?��0��COS��� ��LN#���ߥŴ�  ��=������꼰�<�1Z���VA�MYǱ:���᯻[�THET=0�UNK23�#��l�#ȰCB��CB�#Cz�AS�ѯ����#����SB�#��'GTSkZAC�����&���$DU�phg6�j��E�%eQ%a_��x�NEhs1K�t�� y��A}Ŧկ׍�����LCPH����^U��Sߥ ����������!��(Ʀ�V��V�غ ��UV��V��V
�V�UV&�V4�VB�H��@������d�����H
�UH�H&�H4�HB�O��O��Os���O���O��O
�O�O*&�O4�O(�F�Ҫ��	���SPBA?LANCE_J�6�LE��H_}�SP�>!۶^�^��PFULCb�q����K*1�UTO_<�p�uT1T2�	
22N�q2VP�M�a�� i�Z23	qTu`O��1Q�INSEG2�QREV�PGQgDIF�ep)1�U6�1��`OBK�q�j�w2,�VP�qI�L�CHWAR4B�"A�B��u$MEC�H��J��A��vAX��aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ����C1_ɒT �� x $WEgIGH�@�`$��d\#��I�A�PIFvAN�0LAG�B��S�B�:�BBIL�%OD��`�Ps"ST0s"P�:�pt �!N�C!L ��P 
P2�Aɑ  �2��Tx&DEBU҄#L|0�"5�MMY9C59N��$4�`g$D|1 a$0�ېl� ���DO_:0AK!� �<_ �&� �q�A��B$�"� NJS�8_�P�@���"O�p �� %�T7P?Q��TL4F0TICK,�#�T1N0%�3=pB�0N�P� u3�PR\p��A��5��5U0PR�OMP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a��@RU�COD�#F9U�@�&ID_�P�E�82B> G_SUFF�� �#�AXA�2DO�7/�5� �6GR�#��DC�D ��E��E-��DU4� u�_ H_FI�!�9GSORD�! R 236s�HR�A>N0$ZDT�E�`|�!X5�4 *WL_NA�1�0�R�5DEF_I�X�RF �T�5�"�6�$�6�S�5�UFISm�#�m1|Ј�40c�3�T6�44􁆂�"D� ?rfd�#�D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D�S �D�U�D>b�B�c�E�S �Dd�B�&2v2a�C� ʑ�E�R�E�S�C9wwu�H�0P} d�0,a�ТF0W�h�u�c� ��TE�qY4� }�!LOMB_�r��w0s"VIS��I�TYs"AۑO�#A�_FRI��~SI,a�n�R�07��0R7�3�#s"W�W��Q��%�_���AEAS{#�B��|�x`WB�8�45�55�6|#ORMULA_I����G�W� h �
>75COEFF_O�1&)��1���Go�{#S� 52CA�� :?L3�!GRm� � � $�`4�v2X�0TM�g��`�e�2�c��3ERIqT�d�TAP�  ��LL�Dp`S��_S�Vkd��$�vAP��.���AP� ��SwETU,cMEAG@��@Πt �!HRL � g� (�  0���l��l��aw��RH�0�a�a}d]�d��B��Ay`Gax`��t[Ѐk@REC[Q:q��1SK_A y��� P_!1_USER����*���VEL�����-�!��IzP� �M�T�1CFG��� � �0]O�NGOREJ �0l���~[�� 4 e�8��"�XYZ<S��� 3� ��_ERRK!� U ѐ�1�@Ac�Ȱ�!�>�B0BUFINDX����p� MORy�� H_ CUȱ�1���dAyQ?�I>Q	$ +�a����� �\�G{�� � $SI�h��@2	��VOv�q�- OBJyE| w�ADJUF2�yĈ�AY�����D��OUKP����AMR=�T��-���X2DIR����X8f�1  DYNt�0�-�T� ��R��0� ~���OPWOR��� �,B0SY�SBU����SOP�o���z�Uy�XP�`K���PA�q��Ӭ���OP�@U����}�"1��IMA�G۱_ �п"IM�.���IN������RGOVRD"ё�	���P����  >gplcC��L�`BŰ?l�PMC_E�P�1EN��Mr�1212�R�"�SL| ��� ��R OVSL=S��rDEX\a`��2�:�_"���P#����P������2�C� �P>���#�_Z�ERl���:����� @��:��O�@R	Iy��
[�g@e����s�P�PL���  $FREEY�EEU�~�Z��L����T�� ATU9Sk�,1C_T�����B������p�Vc18��P��� Dc1������LQ����MQ��ۡL�XE��x�5I�P�W�` ��UP��H`&aPX;@���43�� �PG�Y��g�$SUB����q���JMP�WAIT~ ���L�OW���1wē CV!F_A�0��R�Z��CC �R$��28IGNR_PL��/DBTB� P*a�#BW@.t�U�0-�IG��!@I�TNLN,�RBѡb�yN!@��PEED~ >��HADOW� ��t���E������PwSPD��� L_ �A�нP���	#UN�q � �RP (�L�YwPa����PH�_PK���b�RETRIE��x������� H�0NFI���� ���V �$ 2}�d�DBGLV<?LOGSIZz�baKKTU���$D�n�_TXV�EM�!Cڡ��� �-R�#�r>��CHECKz��(��L���ϰq)ҹL��NPA�`T�J"����)1P����
�AR�"�BC =Sa��O�@����ATT S�u䡳&� w�^a�3�-#UX^�4�PL��@Z�� $d��qS�WITCH�h�W���AS��f�3L�LB��� �$BA�Dvc��BCAMi��6I��(@#J5��N�UB6[F
A_KNOWK3qB"ЍU��AD+Hc� D���IPAYLOAq�9p�C_���GrѼG�Z�CLqAj��PL�CL_6� !@4��BOA?�T7�VFYCӐ�Jp��D��I�HRՐ�G�TBd��6�J��zQ_J�A: �B�AND���`�T�BQ�q��PL@?AL_ ��0 P=�TAe��pC��D�C�E���J3�P�V�{ T�PDCK^��)b��COM�_AL3PH�ScBE<�߁��_�\�X�x\� �� ���OD_�1�J2�DDM�AR�<�h�e�f�cQ�TI�A4�i5�i6��MOM(��c�c�c�c�cV�B� AD�cv�c\v�cPUBP�R�d�<u�c<u�b}"�1���� L$PI$� �pc��G�y��I�yI�{I�{I�s�`�A ���v��v�J�bp��a��HIG�3 ���0���5Ѐ0�f�?�5N�5�SAMPD Ƣ�0���8�;@�S ��с 6���1���� ���` ���`1�K�P��`腽P2�H��IN1��P ��8�T�/��:�z�Q��z���GAMM&�S|��$GET�d����D^d>�
$�P�IBR��I��$HI��_���1���E=��A�9�*�LW�W�N�9�{�*�Zb����QCdCHKh0�j�ݠnI_�� M�JļRoh�Q ��s�J�-v��S ý$�X 1�N�I��RCH_D�$RN���^�LE@��i�p�Zh8�ţ_MSWFL/M�P7SCR�75�Ҽ ��3�"Ķ�6��`��`ع�紙��0SV���P'������G�RO�g�S_SA�=AH�=ńNO^`C i�_d=��no�O�O �x�ʚ��p�B�u�ȐcDO�A��!�ں �*�t�:�Z1f�;�7լ���C etMmu�o � �YL�snQ ��� ���"��<s�	�����nQ�8��<3M_Wl���A��\p��(�o�MC ��P���Q���ȇ�hpM.�pr� !��!��$�WM��ANGL�!�AM�6d K�=dK�DdK��TT7�ANk@��3�#�PXC 	OEc�QZ��hp	nt�� ���OM� ��ϑϣϵ����`� �c�Z0���hp^a_�2� |a�J��i ���c���cJ��j������jA�{ �{����{ �@{�P�1�P�MON_QU�� �� 860QCO�U��QTHxH�O��B HYS�0ESPBB UE- 3�f0]O�4�  c P��^�RUN_TOʹ�gpO��� �P�@��IND9E�#_PGRA���0���2��NE_NO���ITf��o INFO��a"��ژ��H�OI� =(*�SLEQ!�*0�*�Q OS��l4�� 460ENA�By� PTION��3��r��^GC]F�!� @60J�,�Q���R�d!���u�PEDITN�� �� ��KAQj"� �E(�NU'�(AUTY�%CO�PYAQ�2,�qe�M��N< @+��PRU�Tm� C"N�OU��2$G��$
�R�GADJ��u2X_��IX����&���&W�(P�(~��&9�� z
�N�P_CYCy�{w�RGNSc9�{�s�LGO£��NYQ_FREQ�SrW@��X1�4�L��@�2P0�!�c@�"�CcRE��MàIF�q��NA��%�4_}Gf�STATU~�<f��MAIL��|CyIq�=LAST�1�a*4ELEMg�� ��QrFEASIt;�ւΰ��B"� F�AF����I� ���O2�E u�vBAB$��PE� =�VA�FzQ�I��TqU[��R���S�FRMS_TRpC�Qc��C��Z�
��1�D � ,2ns�؆�	MB 2� `���N�3V�R 2WR*���шR^W�wNj�DOU�^�N��,2PR`�h�1G�RID��BAR�S!�TYuBOT�Op�� |_"�4!� �R�TO��d�� � ����P�OR�c~vbSReV�0)"dfDI[�T�`;aNd�pXg
�XgQ4Vi��Xg6Vi7ViI8:a�Fʒg�z ?$VALU�C0��3D1@(1F05��C !pf���S�1�-ȆAN/��b�1R��]11ATOTALX����=sPWE3I�Q>StREGENQzfr��X�H�]5	v( cTR�CS�Qq_S3��wfp�V�!��r��BE�3�PG0B�( nsV_H�PDA(��p�S_Ya���i6�S��AR(�2� }�"IG_SE�3ȿpb�5_� �tC_��V$CMPl��D�Ep�G���IšZ�~�X�
�% Fm�HA{NC.� p Q�r�2���INT�9`cq�F���MAsSK�3�@OVRMP �PD�1-��W� ��aХT�l�_RF|�{�V�PSLGP�
g�9�j5��,��;pDpS���4��1U���|�TE���`G���`k���J^�<Y�y3IL_Mx4�s��p��TQ( ����@����V.�C<�P�_ �R�F�M]�V1V\�V1j�2y�2j�U3y�3j�4y�4j� ��p۲������ܲ;IN�VIB8�6��#��*�2&�22�3*&�32�4&�42���6�|�J�  �T ?$MC_FK `� �L>�J�х1p�Mj�Iу��zS ���1���KEEP�_HNADD��!H鴓@�C��0	��Q����
�O!�v ঱�p
�և
�REM!�	�Cq�RF�]�b��U�4e	�HPWD�  �SBM����PCOLLAB�*�p��/q�2I�T/0��""NO1�F�CALp⎵��� �, �FLv�A$�SYN���M��C�k��RpUP_DL�Y��zDELAh9�Dq�2Y AD(���(0QSKIPNO�� �`� O��cNT����c�P_�  ��׾ ��cp���q�� ���o`��|`�ډ`��@�`�ڣ`�ڰ`��9�!O�J2R0  �lX�@TR3H��1AH��� �H���$ RD�Cq��� � R"�R, 5��R�1��8E��5TRGE�_C��RFLG"���9W�5TSPC�1�UM_H��2TH�2N}Q�;� o1� y�ED�Q>02 � D� ˈ<��@2_PC3W��S���1Y0L10_�Cw2$C+��� � $\� U@ ��V7�����0� �� c�\����� r@d��C�Q,��7���DZ Gs�RUVL1b[�1h���10]�_DS�������PK ;11�� lڰ�0���q��AT?��$ �Q[7�� ��K 5Tx���HOME�S *�c2h�n������]�`3h���!3EW `4h�h@z�����5h���	//-/?/W6h�b/t/�/�/�/��/ ���!7h��/�/??'?9?�8h�\?n?�?�?�?�?� _S����  �Aa{p��3��+�_�Ed� T0=�nD4vnCIO䑎I�I@`�O��_OP��E�C.rfBXPOW=E	�� X@��f��$$C�d�S����_��5�3�3� �@�sSI��GP�0�QIRTU�AL�O
QAAVM_WRK 2 7U� ?0  �5Qn_rzXk_�] �\A	�P�]�_3�8P��_�_�Ve�\#m/o�Q`5ojo|o�dHPBS��� 1Y� <Xo�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯz�bC$�AXLM�@tiAQ��c  d��IN����PRE�
�E�J�-�_U�P��[�7QHPIO�CNV_�� �	�Pr�US>��g�c{IO)�V 1U[P $E`��Qս9lҿ8P?��i@��� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o��o�m�LARMRECOV a���-���LMDG ���ɰ�LM?_IF ��� ை����zv����%�6�, 
 6�_��r漅�������̍$w���׏���8�J�\�n����NGTOL  a�� 	 A   ���ț�PPINFoO ={ <v�����1��   I�3�a�"rP���t��� �����ί���>�o����j�|������� Ŀֿ�����0�B��PzPPLICAT�ION ?����J��Handling�Tool �� �
V9.30P/�04ǐM�
88g340�å�F0����202�ťʚϬ�7DF3��M̎��NoneM�F{RAM� 6���Z�_ACTIVE��b  sï�  ~p�UTOMODz��A���m�CHGAoPONL�� ���OUPLED 1ey� �������g�CUREQ �1	e{  T�
��	p��w����#r���e�HN���{�HTTHKY��
$r��\[�m���� O�	�'�-�?�Q�c�u� ������������ #);M_q�� ����% 7I[m��� /���/!/3/E/ W/i/{/�/�/�/?�/ �/�/??/?A?S?e? w?�?�?�?O�?�?�? OO+O=OOOaOsO�O �O�O_�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_oo#o5o GoYoko}o�o�o�o�o �o�o1CU gy������ �	��-�?�Q�c���1�TO��|�p�DO_CLEAN��|n��NM  �� �B�T�f�x����%�DSPDRY�R��m�HI���@ /�����,�>�P�b��t���������ίj�MAXa�ۄ��������Xۄ������p�PL�UGG��܇�ӌ�P�RC��B� ���ׯF�OK���ȔSEGF��K������ �.�����,�>�v���LAPӟ澨�� �϶����������"��4�F�X�j߯�TOT�AL�7���USE+NUӰ�� �������1�RGDISPWMMC����C��&��@@Ȓ��Oѐ������_STRI�NG 1
��
��M��Sl��
A�_ITEM1K�  nl�g�y�� �����������	�� -�?�Q�c�u����������I/O S�IGNALE��Tryout M�odeL�Inp���Simulat{edP�OutOVERRА� = 100O�In cycl�P�Prog A�borP���S�tatusN�	H�eartbeat�J�MH Fauyl��Aler�	 ������*8<N` ׃G� ׁY�c����� ////A/S/e/w/�/��/�/�/�/�/�/wWOR��G�-1�?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO8�O�O�NPOE� �@E;�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo�BDEV�Nu`�Obo�o �o�o�o�o�o, >Pbt��������PALT ��E?�A�S�e�w� ��������я���� �+�=�O�a�s����GRI�G뽑1��� ���	��-�?�Q�c� u���������ϯ�� ��)�����R�a� ՟;���������ѿ� ����+�=�O�a�s���ϗϩϻ���O�PREG��y���-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_��q����$ARG_�-0D ?	������� � 	$��	+[��]����������SBN_CONGFIG���� ��CII_S?AVE  ��)����TCELLSETUP ���%  OME_I�O����%MOV�_Hn�����REP�d�����UTOBA�CKY���#��FRA:\�� �����)�'`l ���&� 7"�� 24/0�6{  09:35:24�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� ,,		�����O�G�O __#_%_7_q_[_�_ _�_�_�_�_�_�_%o����D�@TSK � �M&,O��UP3DT�@EGd�`�F�XWZD_ENB8ED��fSTADE��ܖe��XIS�UNOT 2��&�(��� 	 0|�} Z�0&�? �<_ �/� K��pp�T<�bp�p�8t�}V��)q{|��t�� B=|�o���;9Յ�!{D�x�Q\��gMETc�2Lf�E� P qA|h�iA��A��B-��B��B�y��}?y�J�?��?:��&@5�W?U��s@���}S�CRDCFG 1��� ��z�����ԏ�����Q=���H�Z� l�~�����	�Ɵ-�� ��� �2�D���域���GR�`�`�O���0kNA����	��n��_EDC@1n��� 
 �%-�0EDT-q����L%�p��"���-������������^��  ����2����*�R�bB���*� q���ϧ���3bϮ� @Ͻϯd?�����=�O���sϏ�4.ߞ�{��� ��W���	�߱�?ߏ�5��j�G����#�� ����}�6��6� �Z�����Z����I��7�����&��΀��&m������8^ҿ����	͇� 9K�o��9*�w��	�S��;��CR����B/ T//�/��w//���РNO_DEL�����GE_UNU�SE���IGAL�LOW 1���2p(*SYS�TEM*�s	$SERV_GR�;�B0�@REGK5$8m3�|B0NUMp:�3��=PMU� �u�LAY�p�|?PMPALD@�5�CYC10�.�>x�0�>CULSU�?0�=�2�AM3LOWD�BOXORIt5C�UR_D@�=PM�CNV�6D@1�0�>�@T4DLI��`=O_9	*PRO�GRAJ4PG�_MI�>�OPAL(�E_UPB7_B>�$FLUI_RESU�7p_z?�_�T#MRY>h0�,�/�b �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� ��������"�LAL_OUT �1;l���WD_�ABOR�0?d�I�TR_RTN  �����g�NONgSTOǠ�� 8�CE_RIA_IL0��ۀ��ŀFCFG ��x۔��_LIMY2�2ګ �  �� 	i�J��<�e�g��5��  9��������
����u��PAQPGP ;1�����Q�c�u�4�CK0����+C1��9��@���P�C��CV��]��d
��l��s��P����C[٤m��v���������� C�j���-���?�Â{HE� ONFI�P�q�G�G_P�@1� �%��������ǿٿ����G�KoPAUSaA1�ۃ �B�W��E� ��iϓϹϟ������� ���#�I�/�m��e�����M��NFO �1"��� �7��ߖ��C w��Bb?	�;���8����,,�MA�@�� �ģ�C�Tp���1VC3�����"��3��h3�E�ŀO����c�COLLECT_�"�[�����EN�@��y���k�N[DE��"�3��"1234567890��\1��H ��֕H&��)M� r�\,L�^���]+���� ��������C 2 �Vhz���� ��
c.@R �v���������� ����I�O !���q����u/�/�/�/C'TR��2"'-(׀^)
��.R�#R-�*W�^ 9_MOR�$� �;�l5��l9�?r?��?�?�?�;E2��%JS=,W�?@�@��CR׀K)DցC�R��&u�XOWAWBC4 � A&��׀x׀}A"@Cz  B�@�CG�B8��AC � %��׀ց:�d�43 <#�
�E���I�O�C=A�I��'GM?�C�(�S=���Qd=AT_D�EFPROG ��;%�/m_APIN�USE�V�ۅ�TK�EY_TBL  �s�ہ���	
��� !"#$�%&'()*+,�-./�:;<=�>?@ABCDPG�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������Ga��͓���������������������������������耇����������������������!�PLC�K�\���P�PSTA�n��T_AUTO_�DO��NFsIN�D���n��R_T1wT2N����5�ŀTRLCPLET�E���z_SCR�EEN �_kcscÂU���MMENU 1)O� <�[_#�q� �,�a���>�d���t� ��ӏ����	����� Q�(�:���^�p����� ��̟�ܟ�;��$� q�H�Z���������� Ưد%����4�m�D� V���z���ٿ��¿� !���
�W�.�@ύ�d� vϜ��ϬϾ������ A��*�P߉�`�r߿� �ߨ��������=�� &�s�J�\������������'�,�p_M�ANUAL�EqD�B
12�v�iDBG�_ERRLIP*�{h! 0��������g�NUMLI�M�s:QOE�@DB�PXWORK 1+�{��>Pbt|��-DBTB_�qG ,��kC3!VD�!DB_AWA�Yo�h!GCP �OB=��A�_AL���o�k�Y�p�uO@�`�_�� 1-�+@
-k-6[���_M+pIS�`�@|"@�ONTIM�w��OD��&
��U;MOTNEN�D�_:RECOR�D 13�{ �<�[CG�O�f!T/ [K��/�/�/�/_(�/ �/f/?�/??Q?c?�/ ?�??�?,?�?�?O O�?;O�?_O�?�O�O �O�O(O�OLO_pO%_ 7_I_[_�O_�O�__ �_�_�_�_l_!o�_,o �_io{o�o�oo�o2o �oVo/A�oe P^�
���R ���=��a�s��� �����*�ߏN��� '���ԏ]�̏������ ��ɟ۟v���n�#����G�Y�k�}���TO�LERENC�B��0� L��g�C�SS_CNSTC�Y 24	�t���.������0� >�P�b�x��������� ο����(�:�ä�DEVICE 25ӫ ��ϟ� ������������/��AߟģHNDGDg 6ӫ� CzT�|.!ơLS 27t�S������������/�U�ŢPARAM 8Gb�A��~��RBT 2:�8�<���{CkA� ·�?  � A��8�.SB���A�?B�  ���a������.��  ����A�A�C�����c�u����C�A�D��k�p�z�A�A��HA�c ��A�	�?(uL�^p���A�Bt�/�D��C��_� 	 A=���ABffA#3�3AҊ���AY�A�Cf��a���A�J��7B]���B��Bf�fBᴠ�33Ca$.@R� (�� ���A����
/ ��//)/;/�/_/ q/�/�/�/�/�/�/�/ <??%?r?I?[?m?? �?�?�?�?�?&O8O� PObOMO�OqO�O�O�O �O�O_�OOL_#_ 5_�_Y_k_�_�_�_�_  o�_�_6oooloCo Uogo�o�o�o�o�o�o  �o	h�O�w �����
��.� 	__I'�1_�q��� �����ˏݏ��� %�r�I�[�������� ��ǟٟ&����\�3� E�W����ȯ���ׯ �"��F�1�j�E�s� ����m�������ѿ� 0���f�=�O�a�s� �ϗ��ϻ������� �'�9�Kߘ�o߁��� ��[����(��L�7� p��m������� ����$�����l�C� U���y�����������  ��	V-?�c u����
�� @+dO�s�� ������*/// `/7/I/[/m//�/�/ �/�/?�/�/?!?3? E?�?i?{?�?�?�?�? �?�?�?FO�jOUOgO �O�O�O�O�O�O__ �'O9OO=_O_�_s_ �_�_�_�_�_�_�_o Po'o9o�o]ooo�o�o �o�o�o�o:# 5��O������ ��$��H�Fz�$�DCSS_SLA�VE ;��}�w��`�?_4D  w����AR_MENU <w� >�؏���� �2�^rǏ\�n��\���SHOW 2}=w� � fr [q����Ə�����@,�>�D�b�t��� �� ��ҟϯ����)� P�M�_�q��������� ˿ݿ���:�7�I� [ς�|Ϧ��ϵ����� ����$�!�3�E�l�f� �ύߟ߱�������� ��/�V�P�z�w�� ������������ @�:�d�a�s������� ����\���*�H�N� K]o������ ��28�GY k}������ "�1/C/U/g/y/ �/��/�/�/��// ?-???Q?c?u?�/�? �?�?�/�??OO)O ;OMO_O�?�O�O�O�? �O�?�O__%_7_I_ pOm__�_�O�_�O�_ �_�_o!o3oZ_Woio {o�_�o�_�o�o�o�o Do-Se�o� �o������.�=�O���CFG >�����q��dMC:\���L%04d.CSIV\��pc�������[A ՃCH݀z�v��w�#�  ���:�J�8�S���JP�j�)����p7�-�n�RC_�OUT ?z������a�_C_�FSI ?�� |��� ��@�;�M�_����� ����Я˯ݯ��� %�7�`�[�m������ ��ǿ�����8�3� E�Wπ�{ύϟ����� �������/�X�S� e�wߠߛ߭߿����� ���0�+�=�O�x�s� ������������ �'�P�K�]�o����� ������������(# 5Gpk}��� �� �HC Ug������ �� //-/?/h/c/ u/�/�/�/�/�/�/�/ ??@?;?M?_?�?�? �?�?�?�?�?�?OO %O7O`O[OmOO�O�O �O�O�O�O�O_8_3_ E_W_�_{_�_�_�_�_ �_�_ooo/oXoSo eowo�o�o�o�o�o�o �o0+=Oxs �������� �'�P�K�]�o����� ������ۏ���(�#� 5�G�p�k�}������� şן �����H�C� U�g���������دӯ ��� ��-�?�h�c� u���������Ͽ��� ��@�;�M�_ψσ� �ϧ����������� %�7�`�[�m�ߨߣ� �����������8�3� E�W��{������� �������/�X�S� e�w������������� ��0+=Oxs ������ 'PK]o�� ������(/#/ 5/G/p/k/}/�/�/�/ �/�/ ?�/??H?C?�U3�$DCS_C�_FSO ?�����1 P [?U?�? �?�?�?�?O
OO.O WOROdOvO�O�O�O�O �O�O�O_/_*_<_N_ w_r_�_�_�_�_�_�_ ooo&oOoJo\ono �o�o�o�o�o�o�o�o '"4Foj|� �������� G�B�T�f��������� ׏ҏ�����,�>� g�b�t���������Ο �����?�:�L�^� ��������ϯʯܯg?_C_RPI~>�? �;�d�_�
�}?.�p�����ݿj>SL�@ ���9�b�]�oρϪ� �Ϸ����������:� 5�G�Y߂�}ߏߡ��� ���������1�Z� U�g�y�������� ����	�2�-�?�Q�z� u�������������
 )RM_q� ������* %7Irm�� ���/�ϛ�,� /W/�/{/�/�/�/�/ �/�/???/?X?S? e?w?�?�?�?�?�?�? �?O0O+O=OOOxOsO �O�O�O�O�O�O__ _'_P_K_]_o_�_�_ �_�_�_�_�_�_(o#o 5oGopoko}o�o�o�o �o�o �oHC Ug��������� ����NOC�ODE @������PRE_CHK B���3�A 3��< �7��������� 	 <����� ?#ۏ%�7��[�m�G� Y�������ٟ�ş� !����W�i�C����� y�ïկˏ������ A�S�-�_���c�u��� ѿ�������=�� )�sυ�_ϩϻϕ��� �����'�9���E�o� I�[ߥ߷ߑ������� ��#����Y�k�E�� ��{��������� ��C�U��=�����w� ��������	����? Q+u�a��� ���);_ qg�Y��S�� ��%/�/[/m/G/ �/�/}/�/�/�/�/? !?�/E?W?1?c?�?� ��?�?o?�?O�?�? AOSO-OwO�OcO�O�O �O�O�O_�O+_=__ I_s_M___�_�_�_�_ �_�?�_'o9oo]ooo Io�o�oo�o�o�o�o #�oGY3E� �{�����o �C�U��y���e��� ��������	��-�?� �K�u�O�a������� ��͟��)��1�_� q��}�������ݯ� ɯ�%���1�[�5�G� ����}�ǿٿ���� ���E�W�1�{ύ�G� u����ϯ������/� A��-�w߉�c߭߿� ����������+�=�� a�s�M���ϑ��� ����'��3�]�7� I�������������� ����GY3}� i�������� C/y�e� ������-/?/ /c/u/O/�/�/�/�/ �/�/�/?)?�?_? q?K?�?�?�?�?�?�? �?O%O�?IO[O5OO �OkO}O�O�O�O�O_ �O3_E_;?-_{_�_'_ �_�_�_�_�_�_�_/o AooeowoQo�o�o�o �o�o�o�o+7 aW_i_��C�� ���'��K�]�7� i���m��ɏۏ���� ���G�!�3�}��� i���ş������ 1�C��g�y�S�e��� �������ѯ�-�� �c�u�O�������Ͽ �ןɿ�)�ÿM�_� 9�kϕ�oρ����Ϸ� �����I�#�5�� ��kߵ��ߡ������ �3�E���Q�{�U�g� ������������/� 	��e�w�Q������� ��������+O a�I����� ��K]7 ��m����� /�5/G/!/k/}/s e/�/�/_/�/�/�/? 1???g?y?S?�?�? �?�?�?�?�?O-OO QOcO=OoO�O�/�/�O �O{O�O_�O_M___ 9_�_�_o_�_�_�_�_ oo�_7oIo#oUoo Yoko�o�o�o�o�o�O �o3Ei{U� �������/� 	�S�e�?�Q������� я㏽����O� a�������q���͟�� �����9�K�%�W� ��[�m���ɯ����� ٯ�5�+�=�k�}�� �����������տ� 1��=�g�A�Sϝϯ� �����Ͽ��������Q�c����$DC�S_SGN C�S����#M��22-JUL�-24 11:3{9 E�06��MN��09������ X�L��ԁ����������Дќ�M��Þ��j�����{�VERSION ���V4.2.1�0�EFLOGI�C 1DS��  	D����X�k�X�z�M�PR�OG_ENB  ���b��Л�UL�SE  ����M�_ACCLIM^�������WRSTJNT��v���w�EMO����ѷ�L��INIT� EZ�O��O�PT_SL ?	�S�1�
 	Rg575�Ӆ�74���6��7��5A��1���2��l���G�h�TO  t���.H�]V?�DEX��d�����FPATH ;A��A\4����HCP_CL?NTID ?+�b� l������IAG_GRP �2JS�� �a[�D��  D�� D�  B�  B��@ff��/B!�@[��W�@��q��B�N��C�-Bz���Bp@e`���mp3m7 7�89012345�6�*�[��  �Ao�mAj�1AdA]��
AW|�AP���AJ-AC/A;�A4H|���@�  A��eA�A3!_A�@�@��B4�� ���t���
�u���ApffAj��yAeK�A_�AY��AS� �MC�AF��A@ �O�+/=/O$O�xc K�w(@�X?�8��@��y��/�/�/�/�/8�;�d�2�5?@~f�f@x1'@q���@kC�@d��D@]��@Vv��6?H?Z?l?~?8s��0l��@e�@^��@W\)�@O��@H�0?�<@7K�@.V��?�?�?�?
O8S�@M00G<@A���@<1@5���@/l�@(�w�@!�0�\NO `OrO�O�Ox'g�L_K� ;_�_�__g_�_�_�_ �_o�_�_�_YokoIo �o�o+o�oX�"� �2�17A�@J>���R
q?�33?Y���r��J7�'Ŭ2q63p4��F>r��LJ@��p�Zr�
=@�@�Q�jqZ��@G Ah�@��@��T= c<���]>*�H>�V>�3�>����J<���<��p�q�x��� ��?� �C�  �<(�U�� 4Vr�33��@
���A@��?R�oD��m R�x���Q��t����Z��Џ��؏�,��i?��7N�>�(�>��@Z�=���J�7�G�v�G�J�B��E�����a��@ǐ@����@��@Q��?L �����I�P���&���'��@�K����A�g�q�PC�  C���Cuy�
���ʯ ?����	��Գ�P4���X��v����*Cz�C�8��D�h�3�_�6C �F� ǿB��ֿ����E��T��� =��2������=�?�^>�&$
�I����CT_CON�FIG K|3���eg���STBF_TTS��
����"�����:��{�MAU��~�MSW_CF���L  �OCoVIEW	�MI�U��㯛߭߿��� �������0�B�T� f�x���������� ����,�>�P�b�t� ������������� ��(:L^p� ����� � 6HZl~�������/��RCB�N��!��F/ {/j/�/�/�/�/�/���SBL_FAUL�T O9*^�1G�PMSK��7��TDIAG P���U����q�UD1: 6789012345q2�q���%P�ϭ?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O ��a6�I'�
�?_��TORECPJ?\:
j4 \_�7_[�?�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�O�O_� _�UMP_OP�TION��>qT�RB���9;uPM�E��.Y_TEM�P  È�33B����p�A�pyt�UNI'��ŏq6�Y�N_BRK Q�t�_�EDITOR� q&qh�r_2PEN�T 1R9) � ,&MAIN� A_bpA_IR�VIS$r5� &?COLOC%�b��&DROP_�DEFE�p_3 SO ]�8�v�2���@�w�1��@�x�S�EM|���B�L�B�ARRA_�pNO� ���&PE�G-�ESTEIR�A:���&PI�CKUP��M�P��p 
Ж�&S�EGU2�/����� �&SUMIRP �����F�ؓF���DA_PRENS�A�E����8� �A�F���1_P�LACE0>�H��&
T�5�4�n���&!ؓ/�����R���/�ǯy�b�4��� ٥�/��>��8�J���%EMGDI_S�TA�u~��q���pN�C_INFO 1ySI��b�����`��Կⷮ���1TI� ��o#�Ϡ�0�d�o}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� Hu� �2�D�R�j�R� x������������ ��,�>�P�b�t��� ����������Z�� #5Ga�k}�� �����1 CUgy���� ����	//-/?/Y c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?��? O%O7OQ/GOmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�?Ooo/o�_ [Oeowo�o�o�o�o�o �o�o+=Oa s������_�_ ��'�9�So]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� K�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�C�5�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ���������!� ;�M�W�i�{���� ����������/�A� S�e�w����������� ����+E�Oa s������� '9K]o� ���1����/ #/=G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? ��?�?	OO5/?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�?�_�_o o-O#oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� �_�_����7oA� S�e�w���������я �����+�=�O�a� s���������ߟ� ��/�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��͟׿����'�1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߫�ſ���� �����;�M�_�q� ������������ �%�7�I�[�m���� ���߯��������)� 3EWi{��� ����/A Sew������� ��/!+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�? �?/��?�?�?�?/ #O5OGOYOkO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�?�_ �_�_�_Oo-o?oQo couo�o�o�o�o�o�o �o);M_q ���_����	o �%�7�I�[�m���� ����Ǐُ����!� 3�E�W�i�{����� ß՟矝���/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߩ� �����������1� C�U�g�y������ ������	��-�?�Q� c�u����߫������� ����);M_q ������� %7I[m�� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?���?�?�? �?�OO+O=OOOaO sO�O�O�O�O�O�O�O __'_9_K_]_o_�? �?�_�_�_�_�?�_o #o5oGoYoko}o�o�o �o�o�o�o�o1 CUgy�_��� ��_�	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� �y�����˟�۟� �%�7�I�[�m���� ����ǯٯ����!��3�E�W�i��� �$�ENETMODE� 1U�_�  ���������»��RRO�R_PROG �%��%�����TABLE  ����Q�c�uσ��SEV_NUM ��  �������_AUTO_?ENB  ̵���ݴ_NO�� V�������  *U���������������+���(�:���F�LTR����HIS�Ð�����_ALMw 1W�� ����̍�+;����� ����0�?�_����  ����²u����TCP_VER� !��!��@�$�EXTLOG_R�EQv������SsIZ����STK��������TOL�  ��Dz~���A ��_BWD�U�*�Z�V�ǲ?�DI�D� X��Z�����[�STEP�l�~�����OP_D�O���FACTO�RY_TUNv�d���DR_GRP s1Y��`�d 	p��.° �*u����RHB ���2 ��� �e9 ���b t�o���� ���J5n�YA���A'��q@9�u��
? J�D�� ȸo��_/�(/(�B�  F!A� � @�33R"�3�3-@UUTn*@�P  /ȷ>u.��>*��<�����-E�� F@� �"�5W�%�-J���NJk�I�'PKHu��IP�sF!���-�?�  ?�/9��<9�8�96C'6<�,5���-��YHv ��� ��"�9d����A�FEAT?URE Z�V��ƱHan�dlingToo�l �5��En�glish Di�ctionary��74D St�0a�rd�6�5Anal?og I/O�7�7�gle Shif�t Outo So�ftware U�pdate%Ima�tic Back�up�9SAground Edit�0~�7Camera�0�F�?CnrRnd�ImXC�Lommo�n calib �UI�C�FnqA�@M�onitor�Kt�r�0Reliab<@�8DHCP�IZ�ata Acqu�is�CYiagn�osOA�1[ocu�ment Vie�we�BWual �Check Sa�fety�A�6ha�nced�F�:�Us�nPFr�@�7xt.� DIO �@fi�RT�Wend�PErEr�@LQR�]�Ws�Y�r�0�P E�:FCTN Menu�P�v S8gTP In�'`facNe�5Gi�gE`nrej@p Mask Exc�P�g�WHT^`Pro�xy SvoT�fi�gh-Spe�PS�ki�D�eJP�Pmm�unicN@ons�hurE`'`_�1ab�connect �2xncr``st#ru�2z>peeQP�JQU�4KAREL Cmd. L�`�ua�husRun-;Ti�PEnvkx(`�el +R@sP@S�/W�7Licen�se�Sn\�PBoo�k(System�)�:MACROs�,�b/Offse�@�uH�P8@_�pM�R�@�BP^Mech/Stop�at.p6R"�ui�RKj�x�P�0�P@)�od@wit#ch��>�EQ.����OptmЏ>��`f�iln\=�gw�uulti-T�`tC�9PCM funHw�F�o3T�R?�f�Re�gi�pr�`I�ri�gPFV����0Num� Selb����P Adju�`���J�tatu��
�iZ��5RDM Rob�ot�0scove��1F�ea7��PFreq Anly�g'Rem`��Qn�7F�>R�Servo�P��~�8SNPX b�rvNSN^`ClifQ<ɮBLibr�3鯢�0 q�����o�ptE`ssag?��4��a -C��;��/I_m>B�MILIBk�E�?P Firm6BU��PEcAcck@sKT�PTX_C�eln����F��1�V�or�qu@imulah�A�A�u��Pa�q�U�j@�Ã&�`ev�.B�.@riP޿�USB port- �@iP�PagP��?R EVNT�ϗ�nexcept�P`��t��ſX�]VC�Ar�b�bf�V2PҦ�h$����SܠSCص�V�SGEk�a�UI~�;Web Pl!� �ާ��Խ`�TeQf�ZDT Appl��d�:�ƺ� �Gri=dV�play�R�WD4�R
�.�:n�EQ�+��r-10iA/�7L*��1Grapghic���5dv�S7DCSJ�ck�q�5�larm Cau�se/��ed�8A�scii�a��LosadnP�Upl,�2�Ol�0�AGu�6N�`���yFyc@�r��0���PV��Jo��m� c�R���c���m�./�����Q�2*u:e�RAJ��P�ٶ4eqiqnL����8NRT����9On�0e He�l�HJ�`oI�alletiz?�H������_�tr�[ROS GEth�q��T@e�װ��!�n�%�2D�tP�kg&Up9g~�(2DV-�3D Tri-jQ:EAưDef.qEBa)pdei���, �bImπF�fЎ�nsp.q=�46�4MB DRAM�Z,#FRO5/@e3ll�<�Mshf!r/"�'c%3@pLƖ,ty@s˒xG��m��.[�� ��BUp���Q�B�=mai�P�߫�]Q����@q6wl!u����^`�xR�?eL� Sup������0�P�`cr��@�R����b䚮�pr1uest�rt~QQ��ߋ�L!�4O��q$�K���l Bui7�n���APLCOO�EV�l%��CGU�OCR�G�O��DR��O
TL�S_��BU/_��K��qN_d�TA�OxVB��_�W�ܑZ���_TC�B�_�V�_�W���WF +o�V�O�W._�W�ņoTEH�o�f�O�gt&�oTEj�xVF�_w�_xVGoTwBTw~o2xVH�xVIA��vL�xVLN�yUMz �bo�f_xVN�xV!P���^xVR&xV!S��܇ʏ��W���v���VGF:�L�P2_h��h�V�h��_g�D��h�FFoh���g�RD�� TUT&��01:�L�2V�L��TBGG��v�ra�in�UI��
%HsMI���pon��m�f�"�F�>&KAREL9� ��TPj��<6 SW�IMESTڢF0O�<5�
"a�X�j��� ����ͿĿֿ���'� �0�]�T�fϓϊϜ� ����������#��,� Y�P�bߏ߆ߘ��߼� ��������(�U�L� ^����������� ����$�Q�H�Z��� ~�������������  MDV�z� �����
 I@Rv��� ���///E/</ N/{/r/�/�/�/�/�/ �/???A?8?J?w? n?�?�?�?�?�?�?O �?O=O4OFOsOjO|O �O�O�O�O�O_�O_ 9_0_B_o_f_x_�_�_ �_�_�_�_�_o5o,o >okoboto�o�o�o�o �o�o�o1(:g ^p������ � �-�$�6�c�Z�l� ��������Ə���� )� �2�_�V�h����� ��������%�� .�[�R�d��������� ������!��*�W� N�`������������ ޿���&�S�J�\� �πϒϤ϶������� ��"�O�F�X߅�|� �ߠ߲��������� �K�B�T��x��� �����������G� >�P�}�t��������� ����C:L yp������ 	 ?6Hul ~�����/� /;/2/D/q/h/z/�/ �/�/�/�/?�/
?7? .?@?m?d?v?�?�?�? �?�?�?�?O3O*O<O iO`OrO�O�O�O�O�O �O�O_/_&_8_e_\_ n_�_�_�_�_�_�_�_ �_+o"o4oaoXojo|o �o�o�o�o�o�o�o' 0]Tfx�� �����#��,� Y�P�b�t��������� ������(�U�L� ^�p����������ܟ ���$�Q�H�Z�l� ~��������د���� �M�D�V�h����  H55�2}���21��R7�8��50��J61�4��ATUPͶ5�45͸6��VCA�M��CRI�UI�Fͷ28	�NREv��52��R63���SCH��DOCV�]�CSU��869zͷ0ضEIOC9��4��R69��ES�ET���J7��R{68��MASK���PRXY!�7��OCO��3帨���̸m3�J6˸53���H2�LCH��OP�LG�0�MHCuR��S{�MCS��0��55ضMDS�W���OP�MP�R�M�@�0̶PCM �R0���ض�ж@�51�51<�0n�PRS��69��FRD�FREQn��MCN��93̶�SNBAE�3�SH�LB��M��M���2�̶HTC�TMI�L����TPA��T7PTX��EL�����8������J95n,�TUT�95�wUEV��UEC��wUFR�VCC���O��VIP�CS�C,�CSG8�r�IWEB�HTTf�R6C�N�CG{IG��IPGS)�RC�DG�H7u7��6ضR85�ƷR66�R7��Rn:�R530�680�I2�q�J��H�6<�E6,�RJح�0�4��6o64\�5�N�VD��R6��R8�4Tg����8�9�0\���J93�91Đ 7+���,�D0:oF�CLI����CMS�� �ST�Y��TO�q���7v�NN�ORS�ֱJ% ��j�OL(E�ND��L��Sf(F;VR��V3D���wPBV,�APL��wAPV�CCG䶷CCR|�CD��C�DL@CSBt�C�SK��CT�CT!BL9��U0,(C��y0L8C��TC �y0�'�TC(7TC��CT1E\��07TEh��0V��TFd8F,(GL8)GI�8H�8I��E@\�87�CTM,(M�8UM@8N�8PHHPL8YRd8(TSd8W�In@VGF�GP2���P2���@�H{7VP�D�HF �VPSGVPR�&VT��YP���VTB7Vs�IHb��VI aH'VK��=VGene���� �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=?�O?a?s?�?  H55hT�1�1�[U�3R78�<50ޭ9J614�9AT�U�T�4545�<6έ9VCA�D�3CR�I,KUI8T�528n-JNRE�:52JwR63�;SCH�9/DOCV�JCU�4�869�;0�:EI�O�TsE4�:R69�JESET�;KJ�7KR68�JMA{SK�9PRXYML]7�:OCO\3�<h�J)P�<3|ZJ6�<�53�JH�\LCH^\ZOPLG�;0�Z�MHCR]ZSkMkCS�<0,[55�:�MDSW}k�[OP��[MPR�Z�@�\0n�:PCMLJR0�k�)P�:)`�[51K5u1|0JPRS[�69|ZFRD<JFwREQ�:MCN�:{93�:SNBA}K^�[SHLB�zM�{t�@ll2�:HTC�:�TMIL�<�JTP�A�JTPTX�EL�z)`�K8�;�0�JwJ95\JTUT�[�95|ZUEVZU�EC\ZUFR<JV�CC��O<jVIP�,�CSC\�CSGtlJ�@I�9WEB�:7HTT�:R6{L���CG{�IG[�IP�GS��RC,�DG��[H77�<6�:R�85�JR66JRu7[R|R53{K68|2�Z�@Jml*,|6|6\JR�\	Pj|4L�6�64���5�kNVDZR6+kR84<���IP,��8��90���KJ9&�\91��̫7[KIP�\JD0�F��CL9I�lKCMS�J9�n�:STY,�TO�:��@�K7�LNN|ZO�RS<jJ��MZZ|O]LK�END�:L��S��FVR�JV3�D,�KKPBV\�A�PL�JAPV�ZC�CG�:CCRjC�D�CDL̚CS�B�JCSK�jCTK�CTB��\���\��C�z���CL�TC�LJ�l�TC��TC�ZCTE�J��|�T�E�J��<�TF��FJ\�G��G��l�Hl��I�z)�l�k�CTM�\�M\�M��Nl�P�,�P��R��;�TSr��W��̚VGF��P2��P2�z ��VPDFLJV�P;�VPR��VT��;� �JVTB��V�KIH�VِM�<��VK,�V{�Gene�8�83EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{?��7�0STD~�4LANG�4 �9�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� ��2�D�V�RBT�6OPTNm�������� Ǐُ����!�3�E� W�i�{�������ß�5DPN�4����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}�x�ߡ߳�ted �4 �8��������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������@��ǯٯ�������*�<�N�`�r���9�9���$FEAT�_ADD ?	��������  	��ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu�����DEMO Z��?   ���} ��'��0�]�T�f� �������������� #��,�Y�P�b����� ������������ (�U�L�^��������� ���ܯ���$�Q� H�Z���~�������� ؿ��� �M�D�V� ��zόϦϰ������� �
��I�@�R��v� �ߢ߬��������� �E�<�N�{�r��� �����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo~o �o�o�o�o�o�o�o! *WN`z�� �������&� S�J�\�v��������� �ڏ���"�O�F� X�r�|�������ߟ֟ ����K�B�T�n� x�������ۯү�� ��G�>�P�j�t��� ����׿ο���� C�:�L�f�pϝϔϦ� ������	� ��?�6� H�b�lߙߐߢ����� ������;�2�D�^� h����������� ��
�7�.�@�Z�d��� �������������� 3*<V`��� �����/& 8R\����� ����+/"/4/N/ X/�/|/�/�/�/�/�/ �/�/'??0?J?T?�? x?�?�?�?�?�?�?�? #OO,OFOPO}OtO�O �O�O�O�O�O�O__ (_B_L_y_p_�_�_�_ �_�_�_�_oo$o>o Houolo~o�o�o�o�o �o�o :Dq hz������ �
��6�@�m�d�v� ������ُЏ��� �2�<�i�`�r����� ��՟̟ޟ���.� 8�e�\�n�������ѯ ȯگ����*�4�a� X�j�������ͿĿֿ ����&�0�]�T�f� �ϊϜ����������� �"�,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/
??A? 8?J?w?n?�?�?�?�? �?�?�?OO=O4OFO sOjO|O�O�O�O�O�O �O__9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿����&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t����������   ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�����y  �x�q��� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p��P����q�p�x ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p���������������$F�EAT_DEMO�IN  ��� �����IND�EX���I�LECOMP �[���B���8 SETU�P2 \B~L�  N w�5_AP2BCK� 1]B	  #�)����%����E �	���5 �Y�f��B ��x/�1/C/� g/��/�/,/�/P/�/ t/�/?�/??�/c?u? ?�?(?�?�?^?�?�? O)O�?MO�?qO O~O �O6O�OZO�O_�O%_ �OI_[_�O__�_�_ D_�_h_�_�_
o3o�_ Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0����ׯQ	� P� 2>� *.VRޯ(���*+�Q���W�{��e��PC������OFR6:��ؾg�����T   �2�����\� ��d�*.F��ϕ�	ó����qo�ߓ�STM� 9���ư%�d��ψ���HU߻�Jש�f�x���GIF�A�L��-����ߑ��JPG ����Lձ�n�����#JS�H�����6����%
JavaS�criptt���C�Se���Kֹ�v� %�Cascadi�ng Style Sheets���j�
ARGNAMOE.DT'��OЁ\;��[�k|(>k DISP*rU�Oп��� �
�TPEINS.X3ML/�:\C�cCustom Toolbar���	PASSWOR�D���FRS:�\�� %Pa�ssword Config/c�Q/ �J/�/���/:/�/�/ p/?�/)?;?�/_?�/ �??$?�?H?�?l?�? O�?7O�?[OmO�?�O  O�O�OVO�OzO_�O �OE_�Oi_�Ob_�_._ �_R_�_�_�_o�_Ao So�_woo�o*o<o�o `o�o�o�o+�oO�o s��8��n ��'���]���� �z���F�ۏj���� ��5�ďY�k������ ��B�T��x����� C�ҟg�������,��� P���������?�ί �u����(���Ͽ^� 󿂿�)ϸ�M�ܿq� ��ϧ�6���Z�l�� ��%ߴ��[����� �ߵ�D���h����� 3���W����ߍ��� @����v����/�A� ��e������*���N� ��r�����=��6 s�&��\� �'�K�o� �4�X��� #/�G/Y/�}//�/ �/B/�/f/�/�/�/1? �/U?�/N?�??�?>? �?�?t?	O�?-O?O�?�cO�?�OO(O�O�F��$FILE_DG�BCK 1]����@��� < �)
S�UMMARY.DyG�OsLMD:�O�;_@Diag� Summary�<_IJ
CONSLOG1__&Q_�_NQ�Console� log�_HK	T�PACCN�_o%�o?oJUTP A�ccountin��_IJFR6:I�PKDMP.ZI	PsowH
�o�oKU[`�Exceptio�n�oyk'PMEMCHECK5o�_*_K��QMemory� DataL�F�Al�)6qRIP�E�_$6�Zs%��q Packe�t L�_�DL�$y�	r�qSTAT����S� %~�rStatusT��	FTP���:����Vw�Qmmen�t TBD؏� �>I)ETHERNE���
q�[��NQEthern��p�Pfigura��oODDCSVRAF̏��ďݟd���� verify �all��{D�.���DIFF՟��͟xb��s��diffd���
q��CHG01 Y�@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ��VTRNDIAG.LS�̿޿s�^q=3� Ope���q� SQnostic�EW �)VD;EV7�DATt�Q�xc�u�g�Vis��?Device�Ϫ�IMG7ºo����y�z�s�Imag�n��UP��ES��~T�FRS:\��� �OQUpdates List ��IJg�FLEXEVENQ�X�j߃�f��F� UIF E�v���B,�s��)
PSRBWLOD.CM��sL�������PPS_RO�BOWEL��GL�o�GRAPHIC�S4Dy�b�t���%4D Gra�phics Fi�leu��AOɿ��rGIG���u�
>YvGigE�ة�~�BN�? )��HADOW������\sShadow Chang���vbQRCMERR�n�\s�� CFG Er�ror�tail�� MA��C?MSGLIB� �"^o� ���T�)�ZD�����/XwZD�6 ad�HPNOTI���
/�/Zu�Notific8��H/��AGUO�/ yO?�O'?P?OOt?? �?�?9?�?]?�?O�? (O�?LO^O�?�OO�O 5O�O�OkO _�O$_6_ �OZ_�O~_�__�_C_ �_�_y_o�_2o�_?o ho�_�oo�o�oQo�o uo
�o@�odv �)�M��� ��<�N��r���� ��7�̏[������&� ��J�ُW������3� ȟڟi�����"�4�ß X��|������A�֯ e�����0���T�f� ���������O��s� �ϩ�>�Ϳb��o� ��'ϼ�K����ρ�� ��:�L���p��ϔߦ� 5���Y���}���$�� H���l�~���1��� ��g���� �2���V� ��z�	�����?���c� ��
��.��Rd�� ���M�q �<�`��� %�I��/� 8/J/�n/��/!/�/ �/W/�/{/?"?�/F? �/j?|??�?/?�?�?��$FILE_F�RSPRT  ����0�����8MDON�LY 1]�5�0� 
 �)M�D:_VDAEX?TP.ZZZ�?�?�_OnK6%N�O Back f�ile 9O�4S�6Pe?�OOO�O�?�O __?>_�Ob_t__�_ '_�_�_]_�_�_o(o �_Lo�_po�_}o�o5o �oYo�o �o$�oH Z�o~��C� g��	�2��V�� z������?�ԏ�u��
���.�@��4VIS�BCKHA&C*�.VDA�����F�R:\Z�ION\�DATA\v�����Vision VD�B��ŏ��� '�5��Y��j���� ��B�ׯ�x����1� ��үg�������X��� P��t���Ϫ�?�ο c�u�ϙ�(Ͻ�L�^� �ς��)���M���q�  ߂ߧ�6���Z���� ��%��I�������:�LUI_CONF�IG ^�5|m��� $ h�F{�5������)�;�I���|xq�s��� ��������a���  $6��Gl~�� �K��� 2 �Vhz���G ���
//./�R/ d/v/�/�/�/C/�/�/ �/??*?�/N?`?r? �?�?�???�?�?�?O O&O�?JO\OnO�O�O )O�O�O�O�O�O_�O 4_F_X_j_|_�_%_�_ �_�_�_�_o�_0oBo Tofoxo�o!o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� �����ʏ܏��� $�6�H�Z�l������ ��Ɵ؟ꟁ�� �2� D�V�h���������¯ ԯ�}�
��.�@�R� d�����������п� y���*�<�N�`��� �ϖϨϺ�����u�� �&�8�J���[߀ߒ� �߶���_������"� 4�F���j�|���� ��[�������0�B� ��f�x���������W� ����,>��b t����O���(:�  �xFS�$FL�UI_DATA �_������uRESULT 2`��� �T��/wizard�/guided/�steps/Expertb��/ /+/=/O/a/s/�/�/��*�Conti�nue with{ G�ance�/ �/�/??(?:?L?^?�p?�?�?�? T-�U��90 �`� �?���9��ps�?0OBOTOfOxO �O�O�O�O�O�O�O�  �_/_A_S_e_w_�_ �_�_�_�_�_�_n�?��?�?�<Frip �Oo�o�o�o�o�o �o�o!3E_i {������� ��/�A�S�o$on��HoAO�TimeUS/DST[� �����+�=�O�a��s������'Enabl�/˟ݟ��� %�7�I�[�m������T�?{�ݯ����Æ24Ώ3�E�W�i� {�������ÿտ翦� ���/�A�S�e�wω� �ϭϿ������ϴ�Ư�د� G��Region�χߙ߽߫� ��������)�;�+�America sou�������������)�;��?�y��#߅�G�Y��ditorL������� #5GYk}��+� Touch P�anel �� (�recommen�)���*�<N`r��U���e�w��������accesd�./@/R/d/ v/�/�/�/�/�/�/Q|�Connect� to Network�/(?:?L?^? p?�?�?�?�?�?�?�?
Y���������!/��Introducts߆O�O�O �O�O�O�O__(_:_ U^_p_�_�_�_�_�_��_�_ oo$o6oHo e�Oeo?O�X_�o �o�o�o'9K ]o��R_��� ���#�5�G�Y�k��}�����h`�ooj }oߏ�o��*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ쯫� ��Ϗ1��X�j�|��� ����Ŀֿ����� 0��A�f�xϊϜϮ� ����������,�>� ��_�!���E��߼��� ������(�:�L�^� p���߸�������  ��$�6�H�Z�l�~� ��O߱�s�������  2DVhz�� ������
. @Rdv���� ����/��'/��� `/r/�/�/�/�/�/�/ �/??&?8?�\?n? �?�?�?�?�?�?�?�? O"O4O�UO/yO�O O?�O�O�O�O�O__ 0_B_T_f_x_�_I?�_ �_�_�_�_oo,o>o Poboto�oEO�OiO�o �o�O(:L^ p�������_  ��$�6�H�Z�l�~� ������Ə؏�o�o�o �/��oV�h�z����� ��ԟ���
��.� �R�d�v��������� Я�����*���� ����C�����̿޿ ���&�8�J�\�n� ��?��϶��������� �"�4�F�X�j�|ߎ� M�_�q��ߕ����� 0�B�T�f�x���� ���������,�>� P�b�t����������� ���߱���%��L^ p�������  $��5Zl~ �������/  /2/��S/w/9�/ �/�/�/�/�/
??.? @?R?d?v?�?�/�?�? �?�?�?OO*O<ONO `OrO�OC/�Og/�O�/ �O__&_8_J_\_n_ �_�_�_�_�_�_�?�_ o"o4oFoXojo|o�o �o�o�o�o�O�o�O �O�oTfx��� ������,��_ P�b�t���������Ώ �����(��oI� m��C�����ʟܟ�  ��$�6�H�Z�l�~� =�����Ưد����  �2�D�V�h�z�9��� ]���ѿ����
��.� @�R�d�vψϚϬϾ� �Ϗ�����*�<�N� `�r߄ߖߨߺ��ߋ� տ����#��J�\�n� ������������� �"���F�X�j�|��� ������������ ������u7�� ����,> Pbt3����� ��//(/:/L/^/ p/�/ASe�/��/  ??$?6?H?Z?l?~? �?�?�?�?��?�?O  O2ODOVOhOzO�O�O �O�O�O�/�/�/_�/ @_R_d_v_�_�_�_�_ �_�_�_oo�?)oNo `oro�o�o�o�o�o�o �o&�OG	_k -_������� �"�4�F�X�j�|�� ����ď֏����� 0�B�T�f�x�7��[ �������,�>� P�b�t���������ί �����(�:�L�^� p���������ʿ��� ���џӿH�Z�l�~� �Ϣϴ����������  �߯D�V�h�zߌߞ� ����������
��ۿ =���a�s�7ߚ��� ��������*�<�N� `�r�1ߖ��������� ��&8J\n -�w�Q������ "4FXj|� �������// 0/B/T/f/x/�/�/�/ �/���/?�>? P?b?t?�?�?�?�?�? �?�?OO�:OLO^O pO�O�O�O�O�O�O�O  __�/�/�/?i_+? �_�_�_�_�_�_�_o  o2oDoVoho'O�o�o �o�o�o�o�o
. @Rdv5_G_Y_� }_����*�<�N� `�r���������yoޏ ����&�8�J�\�n� ��������ȟ��� ��4�F�X�j�|��� ����į֯����ˏ �B�T�f�x������� ��ҿ�����ٟ;� ��_�!��ϘϪϼ��� ������(�:�L�^� p߁ϔߦ߸�������  ��$�6�H�Z�l�+� ��Oϱ�s��������  �2�D�V�h�z����� ����������
. @Rdv���� }�������<N `r������ �//��8/J/\/n/ �/�/�/�/�/�/�/�/ ?�1?�U?g?+/�? �?�?�?�?�?�?OO 0OBOTOfO%/�O�O�O �O�O�O�O__,_>_ P_b_!?k?E?�_�_{? �_�_oo(o:oLo^o po�o�o�o�owO�o�o  $6HZl~ ���s_�_�_�� �_2�D�V�h�z����� ��ԏ���
��o.� @�R�d�v��������� П�������� ]����������̯ޯ ���&�8�J�\�� ��������ȿڿ��� �"�4�F�X�j�)�;� M���q��������� 0�B�T�f�xߊߜ߮� m���������,�>� P�b�t�����{� �ϟ����(�:�L�^� p���������������  ��6HZl~ ������� ��/��S�z�� �����
//./ @/R/d/u�/�/�/�/ �/�/�/??*?<?N? `?�?C�?g�?�? �?OO&O8OJO\OnO �O�O�O�Ou/�O�O�O _"_4_F_X_j_|_�_ �_�_q?�_�?�_�?�_ 0oBoTofoxo�o�o�o �o�o�o�o�O,> Pbt����� ����_%��_I�[� ��������ʏ܏�  ��$�6�H�Z�~� ������Ɵ؟����  �2�D�V��_�9��� ��o�ԯ���
��.� @�R�d�v�������k� п�����*�<�N� `�rτϖϨ�g����� ������&�8�J�\�n� �ߒߤ߶��������� ��"�4�F�X�j�|�� �������������� ����Q��x������� ��������,> P�t����� ��(:L^ �/�A��e����  //$/6/H/Z/l/~/ �/�/a�/�/�/�/?  ?2?D?V?h?z?�?�? �?o���?�O.O @OROdOvO�O�O�O�O �O�O�O�/_*_<_N_ `_r_�_�_�_�_�_�_ �_o�?#o�?Go	Ono �o�o�o�o�o�o�o�o "4FXio|� �������� 0�B�T�ou�7o��[o ��ҏ�����,�>� P�b�t�������iΟ �����(�:�L�^� p�������e�ǯ��� ����$�6�H�Z�l�~� ������ƿؿ�����  �2�D�V�h�zόϞ� ���������Ϸ��ۯ =�O��v߈ߚ߬߾� ��������*�<�N� �r��������� ����&�8�J�	�S� -�w���c��������� "4FXj|� �_����� 0BTfx��[� �������/,/>/ P/b/t/�/�/�/�/�/ �/�/�?(?:?L?^? p?�?�?�?�?�?�?�? ����EO/lO~O �O�O�O�O�O�O�O_  _2_D_?h_z_�_�_ �_�_�_�_�_
oo.o @oRoO#O5O�oYO�o �o�o�o*<N `r��U_��� ���&�8�J�\�n� ������couo�o鏫o �"�4�F�X�j�|��� ����ğ֟蟧��� 0�B�T�f�x������� ��ү������ُ;� ��b�t���������ο ����(�:�L�]� pςϔϦϸ�������  ��$�6�H��i�+� ��O������������  �2�D�V�h�z��� ]���������
��.� @�R�d�v�����Y߻� }����ߣ�*<N `r������ ���&8J\n ��������� /��1/C/j/|/�/ �/�/�/�/�/�/?? 0?B?f?x?�?�?�? �?�?�?�?OO,O>O �G/!/kO�OW/�O�O �O�O__(_:_L_^_ p_�_�_S?�_�_�_�_  oo$o6oHoZolo~o �oOO�OsO�o�o�O  2DVhz�� �����_
��.� @�R�d�v��������� Џ⏡o�o�o�o9��o `�r���������̟ޟ ���&�8��\�n� ��������ȯگ��� �"�4�F���)��� M���Ŀֿ����� 0�B�T�f�xϊ�I��� ����������,�>� P�b�t߆ߘ�W�i�{� �ߟ���(�:�L�^� p���������� ���$�6�H�Z�l�~� �������������� ��/��Vhz�� �����
. @Qdv���� ���//*/</�� ]/�/C�/�/�/�/ �/??&?8?J?\?n? �?�?Q�?�?�?�?�? O"O4OFOXOjO|O�O M/�Oq/�O�/�O__ 0_B_T_f_x_�_�_�_ �_�_�_�?oo,o>o Poboto�o�o�o�o�o �o�O�O%7�_^ p�������  ��$�6��_Z�l�~� ������Ə؏����  �2��o;_���K ��ԟ���
��.� @�R�d�v���G����� Я�����*�<�N� `�r���C���g���ۿ ����&�8�J�\�n� �ϒϤ϶����ϙ��� �"�4�F�X�j�|ߎ� �߲����ߕ�����˿ -��T�f�x���� ����������,��� P�b�t����������� ����(:��� �A�����  $6HZl~ =�������/  /2/D/V/h/z/�/K ]o�/��/
??.? @?R?d?v?�?�?�?�? �?��?OO*O<ONO `OrO�O�O�O�O�O�O �/�O�/#_�/J_\_n_ �_�_�_�_�_�_�_�_ o"o4oE_Xojo|o�o �o�o�o�o�o�o 0�OQ_u7_�� ������,�>� P�b�t���Eo����Ώ �����(�:�L�^� p���A��eǟ���  ��$�6�H�Z�l�~� ������Ưد�����  �2�D�V�h�z����� ��¿Կ�������+� �R�d�vψϚϬϾ� ��������*��N� `�r߄ߖߨߺ����� ����&��/�	�S� }�?Ϥ���������� �"�4�F�X�j�|�;� ������������ 0BTfx7��[� �����,> Pbt����� ���//(/:/L/^/ p/�/�/�/�/�/�� ��!?�H?Z?l?~? �?�?�?�?�?�?�?O  O�DOVOhOzO�O�O �O�O�O�O�O
__._ �/�/?s_5?�_�_�_ �_�_�_oo*o<oNo `oro1O�o�o�o�o�o �o&8J\n �?_Q_c_��_�� �"�4�F�X�j�|��� ����ď�oՏ���� 0�B�T�f�x������� ��ҟ����>� P�b�t���������ί ����(�9�L�^� p���������ʿܿ�  ��$��E��i�+� �Ϣϴ����������  �2�D�V�h�z�9��� ����������
��.� @�R�d�v�5ϗ�Yϻ� }������*�<�N� `�r������������� ��&8J\n ���������� ��FXj|� ������// ��B/T/f/x/�/�/�/ �/�/�/�/??�# �G?q?3�?�?�?�? �?�?OO(O:OLO^O pO//�O�O�O�O�O�O  __$_6_H_Z_l_+? u?O?�_�_�?�_�_o  o2oDoVohozo�o�o �o�o�O�o�o
. @Rdv���� }_�_�_�_��_<�N� `�r���������̏ޏ �����o8�J�\�n� ��������ȟڟ��� �"����g�)��� ����į֯����� 0�B�T�f�%������� ��ҿ�����,�>� P�b�t�3�E�W���{� ������(�:�L�^� p߂ߔߦ߸�w�����  ��$�6�H�Z�l�~� ����������� ��2�D�V�h�z����� ����������
-� @Rdv���� �����9�� ]������� �//&/8/J/\/n/ -�/�/�/�/�/�/�/ ?"?4?F?X?j?)�? M�?qs?�?�?OO 0OBOTOfOxO�O�O�O �O/�O�O__,_>_ P_b_t_�_�_�_�_{? �_�?oo�O:oLo^o po�o�o�o�o�o�o�o  �O6HZl~ �������� �_o�_;�e�'o���� ��ԏ���
��.� @�R�d�#�������� П�����*�<�N� `��i�C�����y�ޯ ���&�8�J�\�n� ��������u�ڿ��� �"�4�F�X�j�|ώ� �ϲ�q�������	�˯ 0�B�T�f�xߊߜ߮� ���������ǿ,�>� P�b�t������� ������������[� ߂�������������  $6HZ�~ �������  2DVh'�9�K� �o����
//./ @/R/d/v/�/�/�/k �/�/�/??*?<?N? `?r?�?�?�?�?y�? ��?�&O8OJO\OnO �O�O�O�O�O�O�O�O _!O4_F_X_j_|_�_ �_�_�_�_�_�_o�? -o�?QoOxo�o�o�o �o�o�o�o,> Pb!_����� ����(�:�L�^� o�Ao��eog�܏�  ��$�6�H�Z�l�~� ������s؟����  �2�D�V�h�z����� ��o�ѯ�����˟.� @�R�d�v��������� п����ş*�<�N� `�rτϖϨϺ����� �������/�Y�� �ߒߤ߶��������� �"�4�F�X��|�� ������������� 0�B�T��]�7߁��� m�������,> Pbt���i�� ��(:L^ p���e�w����� ���$/6/H/Z/l/~/ �/�/�/�/�/�/�/�  ?2?D?V?h?z?�?�? �?�?�?�?�?
O�� �OO/vO�O�O�O�O �O�O�O__*_<_N_ ?r_�_�_�_�_�_�_ �_oo&o8oJo\oO -O?O�ocO�o�o�o�o "4FXj|� �__������ 0�B�T�f�x������� moϏ�o�o�,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ���!��E��l�~� ������ƿؿ����  �2�D�V��zόϞ� ����������
��.� @�R��s�5���Y�[� ��������*�<�N� `�r����g����� ����&�8�J�\�n� ������c��������� ��"4FXj|� �������� 0BTfx��� ����������#/ M/t/�/�/�/�/�/ �/�/??(?:?L? p?�?�?�?�?�?�?�?  OO$O6OHO/Q/+/ uO�Oa/�O�O�O�O_  _2_D_V_h_z_�_�_ ]?�_�_�_�_
oo.o @oRodovo�o�oYOkO }O�O�o�O*<N `r������ ��_�&�8�J�\�n� ��������ȏڏ��� �o�o�oC�j�|��� ����ğ֟����� 0�B��f�x������� ��ү�����,�>��P��!�3������$�FMR2_GRP� 1a���� �C4 w B�[�	 [��߿�ܰE�� �F@ 5W��S�ܰJ��NJ�k�I'PKH�u��IP�sF�!���?�  �W�S�ܰ9�<9��896�C'6<,5����A�  l�Ϲ�BHٳB�հ�����@�33�33S�۴��ܰ/@UUT'�@��8���W�>u.�>*���<����=�[�B=���=�|	<�K�<�q�=�mo����8�x	7�H<8�^6�Hc7��x?� ���������"��F��X���_CFG =b»T Q������X�NO ^º
F0�� ���W�RM_CHKTYP  ��[�ʰ�̰����ROM�_�MIN�[����9����X��SSB�h�c�� ݶf�[�]�����^�TP_DEF_�O�[�ʳ��I�RCOM���$�GENOVRD_�DO.�d���TH�R.� dd��_�ENB�� ��RWAVC��dO�Z�� ���Fs  �G!� GɃ��I�C�I(i J���+���%�q���� �Q�OU��j¼��8����<6�i��C�;]�[�C�  D�+��3@���B���p�.��R SMT���k_	ΰ\��$HoOSTCh�1l¹�[��d�۰ M5C[���/Z�  27.0� =1�/  e�/? ?'?9?G:�/j?|?�?�?�,Z?T3	anonymouy �?�?�	OO-O?N�/ڰRH RK�/�?�O�/�O�O�O �O_V?3_E_W_i_�O &_�?�_�_�_�_�_@O �_dOvOSo�_�Ojo�o �o�o�o_�o+ =`o�_�_���� �o&o8oJoL9��o ]�o��������oɏۏ ����4�j+�Y�k� }��������� � �T�1�C�U�g����� ������ӯ��x�>�� -�?�Q�c�����Ο�� �Ͽ����)�;� ��_�qσϕϧ�ʿ � �����%�7�~��� ��߶ϣ�������� ���Ϻ�3�E�W�i�� ���ϱ���������@� R�d�v�x�J��߉��� ���������+ =`���������:$h!ENT 1=m P!V  7 ?. c&�J�n�� �/�)/�M//q/ 4/�/X/j/�/�/�/�/ ?�/7?�/?m?0?�? T?�?x?�?�?�?O�? 3O�?WOO{O>O�ObO �O�O�O�O�O_�OA_ _e_(_:_�_^_�_�_��_�ZQUICCA0�_�_�_?od1@oo.o�od2�olo~o��o!ROUTE�R�o�o�o/!P�CJOG0!�192.168�.0.10	o�SC�AMPRT�\!�pu1yp��vRT��o��� !S�oftware �Operator? Panel�m�n��NAME �!�
!ROBO��v�S_CFG �1l�	 ��Auto-s�tarted'�FTP2��I�K 2��V�h�z������� ԟ����	���@� R�d�v���	����� ��:���)�;�M�_� &���������˿�p� ��%�7�I�[��"� 4�F�ڿ�������� !�3���W�i�{ߍߟ� ��D���������/� vψϚ�w�ߛ��Ͽ� ��������+�=�O� a�������������� ��8�J�\�n�p�]�� ��������� #5X�k}� ���0/D 1/xU/g/y/�/RH/ �/�/�/�//?�/?? Q?c?u?�?���/ ?�?:/O)O;OMO_O &?�O�O�O�O�O�?pO __%_7_I_[_�?�? �?t_�O�_O�_�_o !o3o�OWoio{o�o�_ �oDo�o�o�o�����_ERR n���-=vPDUSI�Z  �`^�P��Tt>muWRD �?΅�Q�  �guest �f������~��SCDMNGRPw 2o΅Wp���Q�`���fK�L� 	P01.�05 8�Q  � �|��  �;|��  ~z[ ���w����*���Ť�x����[ݏȏ���בPԠ�������)����D�r���؊p"*�Pl�P���Dx���dx�*�����%�_GWROU7�pLyN���	/�o���QU%P��UTu� ��TYàL}?pT�TP_AUTH �1qL{ <!iPendan���o֢!KAREL:*�������KC��ɯۯ���VISION SET�9����P�>� h��f�����������ҿ����X�CTRL rL}O�u���a
��hFF�F9E3-ϝTF�RS:DEFAU�LT��FAN�UC Web Server�ʅ�t� X���t@���1�C��U�g�;tWR_CONFIG s;�� ��=qIDL_CPU_PC����aBȠP�� BH��MIN�܅q��?GNR_IOFq{r��`Rx��NPT_S_IM_DO���STAL_SCR�N� �.�INT�PMODNTOL8Q����RTY0���8�-�\�ENBQ�-����OLNK 1tL{�p�������)�;�M���MAST�E�%���SLAV�E uL|�RA?MCACHEk�c�}O^�O_CFG�������UOC�����CMT_OP���Pz�YCL������_?ASG 1v;��q
 O�r��� ����&8pJ\W�ENUMzs5Py
��IP����RTRY_CN���M�=�zs���Tu ������w���p/��p��P_MEMB?ERS 2x;�l�k $��X"��?��Q'W/i)��RCA_�ACC 2y��  X�b� %;�ҿb6���"?� ���Q�&�#�#�/�!����,�$BUF001� 2z�= b�cu0  u0bUs:4�:4�:4�:4U�:4�:4�:4�:4{�C�P^�:3�^��4��4��4Ǫ�4׊4�4�:3_U�4�4.�4@�4�P�4b�4r:3` �V� @`�4!*�40�4B�4Q�494�`A4`��4��4���4��4��4��4�Z�4�:3azD zDVDaCzDSzDdzD�tzDADaIDaY4aU�zD�zD�zD�zDU�:4:4:4/:4�4b�492$?63:1 @1ERI0ERQ0ERY0ER a0ERi0ERq0ERy0ER �0�1�1:1�1�R�0�R �0�R�0�R�0�R�0�R �0:1�1�R�0�R�0�R �0�R�0�R�0�R�0:1  AAAb@b@b !@b)@bBT8AbA@ bI@bQ@bY@ba@ bi@bq@by@:1�A �b�@�b"d�A�b�@�b �@�b�@�bJd�A�bbT �A�b�@�b�@�b�@�b �@ER�@ERPER	PER�TQ:193-_65GS NrI2WSNrY2gSNri2 wSNry2�S���3�S�r �2�S�r�2�S�r�2�S ���3�S�r�2�S�r�2 �S�r�2c�	Bc� B'c�)B7c�St@C Oc�QB_c�aBoc� qBc���C�c��+��C �c���B�c��S��C�c ���B�c���B�c���B �cNrRsNr�tS'v��2{�4r�}ŋ���<����o�o��2�HIS!2}�� ܷ! 2024-07-22��A��П����`�� o�� m�)�;�M�_�o��X�fn��6-2�7������Ư�ɕr;0����fn#��p"�4�F�}��g��6��~�����ٮo��o���g������\"�}��j���5m��Z�l�~�٬ 7 5�h�j����p������y��cN���1O�L�9�K�]�ܩ/ 9 ɽcP����߸�������mv��0l��#�5﴿�;Z�M 9 ��h�mv{�;M }�����`���!	���� �,�>�P�b�t���i ��,P����������#�;{�b� o�d ,_q�q���������M��c��d >K ��I6HZl Z� ���H�%� %ٰ%/$/6/H/�6�H�~/�/�/�: B�����/�/ ??��(?g?y?�?8�P�"�" a�� �/�?�?�? O�ߑ6O�HOZOH�&  @e�Ac�"C u�o�chO�O�O�O�����O _1_C_U_g_y_�_�_ �_����5p����(Oo$o6oHo6�secro �o�o�o��o�o M�fb�fbce��no [m�%O�� �"4رJ7�I�[��m�[/m/����ǏH� ��> ꂵ�fb��&� �-�?�-???������@��P��B��B> p� ��֒�����OO s�`�r���M��L�e�����u���ԯ� ���O�OS�@�R�d�v����������п�_�RI_CFG 2~�[� H
Cycle Time��Busy�I�dl��minz�S�Upƾ�Read(��DowG�C�{���Count>�	Num �������L�����P�ROG���U��P�)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,1�C�U��g�y�Tä�SDT_�ISOLC  ��Y� ���J2�3_DSP_EN�B  ��T���INC ���L����A   ?�  �=���<#�
|���:�o ��2�D�L�/�l���OB���C��O��ֆ�G�_GROUP 1큦��<�*�����t�?����L�Q'�L�^�p�@/����������\��~�G_IN_AU�TO����POSR�E���KANJI_MASK0��D�RELMON ��[��L�y����@����f�Ã�ǉ��L�-��K�CL_L NUM���G$KEYLO�GGINGD�P�������LANGU�AGE �U���DEFA�ULT ��QLGf�����S��L��xస�8T�H [ �L�'0��L���!��K�L�;��
�*!(UT1:\ J/ L/Y/k/}/ �/�/�/�/�/�/�/$>�(�H?�VLN_D?ISP ���P��&�$�^4OCTOL��Dz����
�1GBOOK ��Ad4V�11�0�� %O!O3OEOWOiKyM0�TËIgF	�5)�����O}���2_B�UFF 2���# �L��U_�2 ��6_M�R_d_�_�_�_ �_�_�_�_�_o3o*o <oNo`o�o�o�o�o��~�ADCS ��� ���L�O��+=�Oa�dIO 2���k +����������� �*�:�L�^�r����� ����ʏ܏���$��6�J�uuER_ITM��d������ǟٟ ����!�3�E�W�i� {�������ïկ���8��7x�SEVD��]t�TYP�����s������)RST�e�eSCRN_F�L 2��}��� ��/�A�S�e�w�F��TP{��b��=NGNAM��E�n�dUPSf0GI���2����_LO{AD��G %��%DROP_�?EITO_3�ϑ��MAXUALRMXb2�@���
K�N��_PR��2  �34�AK�Ci0��qO�=_'X�Ӭ�P 2���; �*V	����
* ���4�� *��'�`�	xN��z� �����������1� C�&�g�R���n����� ������	��?* cFX����� ��;0q \������� /�/I/4/m/X/�/ �/�/�/�/�/�/�/!? ?E?0?i?{?^?�?�? �?�?�?�?�?OOAO�SO6OwObO�OD�DBG*� ��գѢ���O�@_LDXDI�SA����ssMEM�O_AP��E ?=��
 �Ax $_6_H_Z_l_~_�_�_�K�FRQ_CFG� ����CA �w@��S�@<��dA%�\o�_�P�Ґ�����*zZ`/\b **:eb �DXojho�F�o�o�o �o�o�o;�O�ՀdZ�U�y|��z,(9�Mt���1� �B�g�N���r����� ���̏	���?�A�?ISC 1���K` ��O�����O���O�֟����K�]�_MS�TR �3��S_CD 1�]�� l��{�����دï կ���2��V�A�z� e�������Կ����� ��@�+�=�v�aϚ� �Ͼϩ��������� <�'�`�K߄�oߨߓ� ���������&��J� 5�Z��k������ ��������F�1�j� U���y����������� ��0T?x�MK�Q�,��Q�$MLTARM�R��?g� �~s�@���@METsPU�@l��4��NDSP_ADC�OL�@!CMNmT7 *FNS|W(FSTLIxi%� �,�����Q��*POSC�F�bPRPMlV�ST51�,�w 4�R#�
g! |qg%w/�'c/�/�/�/ �/�/�/?�/?G?)? ;?}?_?q?�?�?�?�?��1*SING_C�HK  {$M7ODA�S�e����#EDEV 	��J	MC:WLHOSIZE�Ml �#ETASK %�J�%$123456�789 �O�E!GT�RIG 1�,� l�Eo#_�y_S_��}�FYP�A�u9D�"CEM_INF �1�?k`)�AT&FV0E0�X_�])�QE0V�1&A3&B1&�D2&S0&C1�S0=�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_ �_o�3o��o�� �o��"�4��X� ��ASe֏�� �C�0���f�!��� q�����s�䟗����� ͏>��b���s���K� ��w���ٯ�ɟ۟ L����#�����Y�ʿ ����$�߿H�/� l�~�1���U�g�y��� �ϯ� �2�i�V�	�z��5ߋ߰ߗ���PONIwTOR�G ?kK�   	EX�EC1o�2�3��4�5��@�7*�8�9o�� ����(��4��@� ��L��X��d��p⨂�|��2��2��2���2��2��2��2���2��2��2��3ʉ�3��3(�#AR_�GRP_SV 1ݛ�[ (�1@3�>�?|�/�Q���6 `��@?Q�>��zRM�A�_DsҔN��ION�_DB-@�1Ml/  �l CFH"�?+�qGG��N� BL"FI-u�d1}E���)P�L_NAME �!�E� �!D�efault P�ersonali�ty (from� FD)b*RR�2�� 1�L��XL�p�X  d�-?Qc u������� //)/;/M/_/q/�/�/�/f2)�/�/�/ ??,?>?P?b?t?f<�/�?�?�?�?�?�? 
OO.O@OROdOc	�6��?�N
�O�OfP �O�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_�O�O2oDoVohozo �o�o�o�o�o�o�o
 .@o!ov�� �������*��<�N�`�r����� �Fs  GT�G�Me��x �ÏՍfd����� ��(�6������
 ��m�~�h�����  ������ğ֟�����@:���
�]�m�f���	`������į��:�oAb	������ A�   /���P����r����� ��^�˿ݿȿ��%�:�R�� 1��	X ���, � ���� a� @D�  t�?�z�`�><|�fA/��t�{	ު�;�	l��	 ��x�J������ �� ��<�@���� ���·�K�K� ��K=*�J����J���J9��
�ԏC����t�@{S�\��(Ehє��.���I����>����T;f�ґ��$��3��´  �@��>�Թ�$��  >�����{�Uf��x`���� �
��������� �  _{  @T����_�  �  �l��ϊ�-�	'� �� ��I� ��  �<�+�:��È��È=̣����0Ӂ��N �~[��n @� ��f���f�k���x,�av�  '������@2��@��0@�Ш���C���Cb C��\C��������@%������� )�Bb $/�!��L��Dz�o�ߓ~���0��( �� -����0����!���/�����恀?�ff0G�*<� }�qD�1�8����>��Hbp��(�(���P���	������>�?�՚��x���W�<
�6b<߈;����<�ê<�?��<�^��I/2��A�{��fÌ¾,�?fff?_�?y&� T�@�.�"�J<?�\��"N\�5���!��(� |��/z��/j'��[0? ?T???x?c?�?�?�?`�?�?�?5��%F� �?2O�?VO�/wO�)IO��OEHG@ G@�0��G�� G} ଙO�O�O_	_B_-_\f_Q_BL��B[�Aw_[_�_b��_�[�_ ��mO3o�OZo�_~o�ox�o�o���b��PV( @|po	lo- *cU�ߡA���r5eCP�Lo�}?����#���5��W�s��6�Cv�q�CH3� j�t�����q�����|^(�hA� �AL�ffA]��?��$�?��;����u�æ�)��	ff��C��#�
���g\)��"�33C�
������<��؎G�B����L�B�s?����	";��H�ۚG��!�G��WIY�E���C�+��8�I۪I�5��HgMG��3E��RC�j�=x�
�pI����G��fIV=�E<YD�C <�ݟȟ����7�"� [�F��j�������ٯ į���!��E�0�i� T�f�����ÿ���ҿ ����A�,�e�Pω� tϭϘ��ϼ������ +��O�:�s�^߃ߩ� ���߸������ �9� $�6�o�Z��~��� ���������5� �Y� D�}�h�����������@����
C.(�g���/"���<��t��q�3�8����q4�Mgu���q�V�wQ�
4p�+4�]$$dR��v���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/��/�/�/�/  %� �/�/+??O?:?s?/`�_�?�?�?�;�?��?O�? OFO4O�r LO^O�O�O�O�O�O�J  2 Fs�w�GT�V�M��uBO�|r�pp�C��S@�R_�to}_�_hf_�_�|\!�W�Ƀ�_oo(o�z?_���@@�z�D��p�pk1�p�~
 6o�o�o�o �o�o�o);M�_q�ڊsa �����D��$M�R_CABLE �2�� �]��T�LaMa?��PMaLb�p�Z���&P�C�p�!O4>ߔB����!Y�4� �!E�h�\�&��v�l  ���&P�v�wdN��{0��$s8<ca��F�� 6��H�XT��6P� C$��Č��n���	� 'z�"�,����� ��&P���C���=��������� )z��~։��s9��T� ,�>���b�������Ɵ ��Ο3�.��P�(�:�@��^���j��#� �� ����;h�H�Z�l��;h*��** ��sOM ��y����B�"%K�%% 23456�78901ɿ۵ �ƿ���� �� AQ�� �!
�z��not sent� ���W��TESTFECS7ALG� eg;jAQ�d��ga%�
���@���$�r�̹�������� 9UD1�:\mainte�nances.x�mS�.�@�vj��DEFAULT��\�rGRP 2�^��  p� �J��%  �%1s�t mechan�ical che�ck��!���������E��Z��(�:�L�^ﾳ��co�ntroller �Ԍ��߰��D���`�� ��$���M��L��""8b���v��B������������/�C}�a�6�����dv���s�C���ge��. battery�&��E	S(:L^pܿ	|�duiz�ab;let  D�а�R����/"/4/���grgeas��'f�r#!-� |!�/�E��/��/�/�/�/��
�oai,�g/y/�/�/@t?�?�?�?�?���
$�XֈW��1<X�AO�E
c?8OJO\OnO��O�t��?O���'O�O_ _2_D_��OverhauE�6�L��R xXЌQ�_���O�_�_�_�_oX�$�_0o����_o �_�o�o�o�o�oo �o?oQocoJ\n ���o�)� �"�4�F���|�� k��ď֏����[� 0�B���f��������� ��ҟ!���E�W�,�{� P�b�t�����矼�� ��A��(�:�L�^� ����ѯ㯸��ܿ�  ��$�s�Hϗ���~� Ϳ�ϴ�������9�� ]�o�Dߓ�h�zߌߞ� ������#�5�G���.� @�R�d�v��ߚ����� �������*�y��� `���O���������� ��?�&u�J��n �����); _4FXj|� ���%�// 0/B/�f/���/� �/�/�/�/?W/,?{/ �/b?�/�?�?�?�?�? ?�?A?S?(Ow?LO^O pO�O�O�?�OOO+O �O_$_6_H_Z_�O~_ �O�O�O�_�_�_�_o8 o�P�R	 T"oOo aoso�_�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
���  ��Q?� ; @�a �oW� i�{��fC�����̟aXw*�** �Q �V��� �2�D��h�8z��������_�S ������կ7�I� [�����ɯ/���ǿٿ #���!�3�}����� {ύϟ��s������� C�U�g��S�e�w�9�@�߭߿�	�߉e�a��$MR_HIS�T 2��U��� 
 \jR$ 2�34567890�1*�2����)�9 c_���R��a_���� �����=�O�a��*� x�����r����� ��9��]o&�J �����#� G�k}4��d��SKCFMAP � �U������`��ONREL  �����лEXC/FENB'
���!FNC$/$JO�GOVLIM'd��m �KEY'zp%y%_PAN(��"�"�RUN`,��+SFSPDTY�PD(%�SIGN|/$T1MOTb/�!�_CE_G�RP 1��U �"�:`��n?�c[?�? �؆?�?~?�?�?�?!O �?EO�?:O{O2O�O�O hO�O�O�O_�O/_�O (_e__�_�_�_�_v_��_�_�_o�׻QZ_EDIT4��#�TCOM_CFG 1��'%to�o��o 
Ua_ARC�_!"��O)T_M�N_MODE6=�Lj_SPL�o2&UAP_CPL�o�3$NOCHECK� ?� � Rdv��� ������*�<��N�`��NO_WA�IT_L 7Jg50N�T]a���UZ޲�_ERR?12���ф��	��-�����R�d����`O�����| %��
aB�����o����C�������,V9<� �� ?�Uϟ�j����قPARAuMႳ��N��oR�=��o��� = e������گ� ȯ��"�4��X�j�F�<�蜿��A�ҿ�"?ODRDSP�c6�/(OFFSET_�CAR@`�o�DI�S��S_A�`A�RK7KiOPEN_FILE4�1�a�Kf�`OPTION�_IO�/�!��M_�PRG %�%c$*����h�WOT�[�E7O��и�Z��  ��� �Z"�÷"�	� �V"�Z����RG_DSBOL  ��ˊ����RIENTT5O ZC����A �U�`IM_ED���O��V�?LCT ���Gb�ԛa�Zd��_P�EX�`7�*�RAT��g d/%*��UOP ���{��������������$�PAL�������_?POS_CHU�7�����2>3�L��XL�p��$�ÿU�g�y����� ����������	- ?Qcu����Y2C���"4 FXj|��� ��� //$/6/H/ Z/l/~/�Y���.��/�/ςP�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO�/�/ LO^OpO�O�O�O�O�O �O�O __$_6_H_Z_ )O;O�_�_�_�_�_�_ �_o o2oDoVohozo`�o�o�_<���o�m ���~B Pw�m�m���~�jw8��w����� �2�T��p��w���H��t	`���̏ޏ��:�o����� �|2��pA�  I� �j�`�������� �џ���@��#��)�Or�1��_�� 8���, �\Ԡ��� @D�  ��?����~�?� ���!D�������G�  �;�	l��	 ��xJ�젌����� �+<� ���%�	��2�H(��H3k�7HSM5G�2�2G���GNɁ3%�R��oR�d�2�C%f��a��{�ׄ���|��/��3��¸��4��>���К������3�A�q½{{q�!ª��ֱ� "�(«�=�2�ܤ��� ��{ � @�Њ���  ��Њ�2����.�	'� � ���I� � � �V�,�=�������˖ß��� � �y��n �@"��]�<߼+��ȅ���-�N�Д�  �'�Ь�w�ӰC��C��\C߰��Ϲ�x�ߤ!���@�4�I��/��2�~�B��@B�I�;�)�j客z+����쿱����������( �� -��#������&�!�]�9��  q�?�ffaH�Z���� ��������8� ����>�|P��}�	(� ��P�������\�?��� x�� ���<
6b<�߈;܍�<��ê<���<G�^�*�gv�A)�ƙ�脣��F�?f7ff?}�?&� ���@�.��J<�?�\��N\� �)���������� �ޤy�N9r] �������/ &/�J/5/n/�	�g/�/c(G@ G�@0i�G�� G}���/??<?'?`?�K?�?o?BLi�B��A�?y?�?|��?K �?ů�/QO�/xO�?�O�O�O�Om��b��n�t @|�O'_�O@K_6_H_�_lS��A��RS�i�Cn_�_j_0O�]?��ooAol,o¹�Wi���To3C���`CHQo>J�d�`a�a@I�ܚ>(hA� ��ALffA]���?�$�?����ź°u�æ��)�	ff��?C�#�
�op�g\)��33C��
�����<���nG�B����L�B��s�����	0źH�ۚG���!G��WI�YE���C��+�½I۪�I�5�HgM�G�3E��R�C�j=�~
�p�I���G��f�IV=�E<YD�#Zo���
� �U�@�y�d������� ��я�����?�*� c�N���r�������� ̟��)��9�_�J� ��n�����˯���گ �%��I�4�m�X��� |���ǿ���ֿ��� 3��W�B�Tύ�xϱ� ����������	�/�� S�>�w�bߛ߆߿ߪ� ��������=�(�a�:L�(q��)�����Z��x����a3�8���<���a4Mgu�����a�VwQ�(�4p�+4�]B� B���p����������U%PbP���QO%�x�1[FjR��������  C���I4m X�8
O������.//>/d/R/�Rj/|/�/�/�/��/�/:  2 {Fs�gGT�&6�M�eBmp�R�P�aC��3@�_p?�?@�?�?�?�?�=�S��OO)O;OMO�c?̯��@@�j�R�`�`�1�`�^
 TO�O�O�O�O �O_#_5_G_Y_k_}_p�_�_�j�A ������D��$PA�RAM_MENU� ?B���  DEFPULSE{�	WAITTM�OUTkRCV�o SHEL�L_WRK.$CUR_STYL`;DlOPTZ1Zo�PTBooibC?oR?_DECSN`�� �l�o�o�o& OJ\n�������QSSREL_�ID  >�
1���uUSE_PRO/G %�Z%�@��sCCR` �
1�S�S�_HOST �!�Z!X���M�T  _���x������>L�_TIMEb ��h��PGDEBU�G�p�[�sGINP?_FLMSK�E�qT� V�G�PGAr�e 5��?��CHS�^D�TYPE�\�0��
�3�.�@�R� {�v�����ï��Я� ���*�S�N�`�r� ���������޿�� +�&�8�J�s�nπϒ����G�WORD ?�	�[
 	PyR2��MAI�`ΓSU�a��TE�Ԁ���	Sd�CCOL��C߸�L�� C�~�h�d�*�TRACECToL 1�B��Q� ��m n�'��0�ށ�DT� Q�B��М�D � ��q����������1�@�@�@���@�@� �U �	������U�����&��.�U��������U�&��.��6��>�U�F�
H�H�H����������� RH� ���������M�������U�����&��.��6��>�U�g�y����G�����������+ �������� ����/�A�S�e�w� ���������������������O��O�O�Ug�X���XXXX��Xf����V��V�V�V��V���V��V��V��V*��V��V�ѐ!�������@����  2DNhz�f ����-�?����? �?�?����������d5 (O:OLO^OpO�O�O�O �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� P�$Or���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~�f������  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o�o�o�o�a�$PG�TRACELEN�  �a  �_��`��f�_UP �����q'pq� p�a_CFG M�u	s�a p�LtLtfqwpqz�  �qu4rD�EFSPD ��?|�ap��`H�_CONFIG s�us �`��`d�t��b ��a�qP�t�q��`���`IN7pTRL' �?}_q8�u��PE�u��w��qLt�qqv�`LI�D8s�?}	v�LL�B 1��y k��B�pB4Ńqv �އ؏	��s << �a?��'���A� o�U�w�������۟���ӟ��#�	�+�Y�v� 񂍯����ï
���������/�u�GRP �1ƪ��a@俼j��hs�aA��
D�� D�@� Cŀ @�٭^�t�q�����q�p���.� ���FȾ´���ʻB� )�	���?�)�c��a�>��>�,���Ϻ��ζ� =49X=H�9��
��� �@�+�d�O���s߬��o߼�����  Dz���`
��8���H� n�Y��}������� ������4��X�C�|����)��
V7.10beta1Xv A�������!�����?!G��>\=y��#��{33A!�ߚ@��͵��8�wA��@� A�s�@Ls���� ��"4FXLsA�pLry�ā���_��@l��@ë33q�`s��k���Anff�a���ھ��)�x�� �ar�T� n�t����	t��KNOW_M  �|uGvz�SV ��z�r�&�� ��>/�/G/�aԤ�y�MM���{ ����	^u (�l+/�/',_t@oXLs�����@���%�"4�.�N�z�MRM��|-T�U�y�c?u;eOADBANFWD~�x�STM�1 1��y�4Ga�rra_B�2Se�m��?~s�;CEo�2��O�7�3�Antena_F?ull @��VO De�qH��^OpO�O�O �O�O�O�O!_ __W_ 6_H_�_l_~_�_�b�7�2�<�!4�_  �#<�_�_N�3�_�_
oo�749oKo]ooo��75�o�o�o�o�76 �o�o�772DVh�78����V�7MA�0��s�wwOVLD  ��{�/a�2PAR?NUM  �;]���u�SCH*� �8�
����ω�3�U�PD��[�ܵ+�wu_CMP_r -��0��'�5C�ER_C;HKQ����1�"e�N�`�RS>0�?G�'_MO�?_��#u�_RES_G�0��{
Ϳ@�3�d�W� ��{��������կ����*�����P� �O��8`l������ �`��ʿϿ��`�	� ��1p)�H�M���p hχό���p�������V 1��5�1�!�@`y�ŒTHR_INR>0/�Z"z�5d:�MASSGߛ Z[�MNF�y�M�ON_QUEUE� ��5�6Ӑ~  U#tNH�U��N������END������EXE�����BE�������OPTIO�������PROGR�AM %��%���߰���TASK�_I,�>�OCFG� ά�]�����D�ATAu#�����Ӑ2�%B�T�f�x� ��5��������������,>P�INFOu#� ����� ����'9 K]o�����@���/lx� �c ;���ȀK_������S&ENB�-�b-&q�&2�/�(G���2�b+ X,�		��=���/��@��P4$��0��99)�N'_E?DIT ���W?|i?��WERFL��-ӱ3RGADJ {�F:A�  �5�?Ӑ�5Wј6��]!�����?�O  Bz�WӐ<1Ӑ�%�%O�8;��5f0!2��7�	H��ml0�,�BP�0��@�0�M�*�@/�B **: �B�O�F�O2��D��A�ЎO�@O	_,X��t%���H�q��O�$_r_0_�_���Q@WA ��>]�_�_�_o�_o �_�_
o�o.o�ojodo vo�o�o�o�o�o�o\ XB<N�r� ���4��0��� &���J���������� �������x�"�t� ^�X�j�䟎���ʟğ ֟P���L�6�0�B��� f���������(�ү$� �����>���z�t� �� Ϫ������l�@�h�R�L�^�DX	����ώ0�� ���t$ :�L��o�
ߓߥ���7PREF ���:�0�0
�5IOORITYX�M6��1MPDSPV�:
B� �UT��C�6OD�UCT��F:��NFOG[@_TG��0��J:?�HIBI�T_DO�8��TO�ENT 1�F;� (!AF_I�NE*�����!�tcp���!�ud��8�!iccm'��N?�XY�3��F<��1)� 0�A�����0����� ������' ] D�h�����$�*>��3��9
BpOTf�3>���2
�B�G/�LC��4��;LFJAB,  ���F!//%/(7/�5�F�Z�w/Љ/�/�/�3&EN�HANCE �2FBAH+d�?�%D;�������Ӓ1�1�PORT_NUM�+��0���1_�CARTRE�@|��q�SKSTA*�ު�SLGS������C�Un?othing?�?�OO�۶0TEMPG �N�"O�E�0�_a_seiban|߅OxߕO�O�O�O �O_�O'__K_6_H_ �_l_�_�_�_�_�_�_ �_#ooGo2okoVo�o zo�o�o�o�o�o�o 1U@e�v� ���������Q�<�u�.IVERS�I	�L��� disable��.GSAVE ��N�	2670H�771|�h��!`�/��9�:� 	^�H4�ϐ����e�� ͟ߟ�����9��D�C-Å_y� 1�
������ő�x���Ǻ�URGE� 1B��r�WFϠ��-��9�W����l:�WRUP_DEL�AY �=n�W�R_HOT %���7��/p��R_NORMALO�V�_�<����SEMI����|����QSKIPo�	�97��xf�=�b�a� sυ�H��ʹ��ø��� �����&��J�\�n� 4�Fߤߒ������߲� ��� �F�X�j�0�� |����������� 0�B�T��x�f����������ãRBTIF��5���CVTMO�U�7�5���D�CRo��� ��T�A�:CC��avC�>��;P>�[a:��_�H�� �c���^��?��S�`kϻ4�HϘ�� <
�6b<߈;����>u.�>*?��<��ǪP0���2DV hz��������,GRDIO_T?YPE  v���/ED� T_CF�G ��-�BHf]�EP)�2��+7 ��B�u �/ �*��/�?�/%?= �/V?�}?�Ϟ?���? �?�?�?�?O
O@O*G l?qO��8O�O�O�O�O �O�O�O�O_<_^Oc_ �O�__�_�_�_�_�_ o�_&oH_Mol_o�o o�o�o�o�o�o�o�o "DoIho*j� ������.3� E��f� ���x����� ���ҏ�*�/�N�� b�P���t�����Ο���ޟ�:�+���R'INOT 2�R��!�1G;� i�{��"�<��8f�0 ��ӫ ������M�;� q�W�������˿��� տ�%��I�7�m�� eϣϑ��ϵ������� !��E�3�i�{�aߟ� ���߱����������A���EFPOS1� 1�!)  x���n#����� ��������/��S� ��w����6�����l� ������=O���� 6���V�z � 9�]�� ��Rd���#/ �G/�k//h/�/</ �/`/�/�/??�/�/ ?g?R?�?&?�?J?�? n?�?	O�?-O�?QO�? uO�O"O4OnO�O�O�O �O_�O;_�O8_q__ �_0_�_T_�_�_�_�_ �_7o"o[o�_oo�o >o�o�oto�o�o!�o EW�o>��� ^�����A�� e� ���$�����Z�l� ����+�ƏO��s� �p���D�͟h�񟌟 �'�ԟ�o�Z��� .���R�ۯv�د��� 5�ЯY���}���*�<� v�׿¿����Ϻ�C��޿@�y��e�2 1�q��-�g�����	� �-���Q���N߇�"� ��F���j��ߎߠ߲� ��M�8�q���0�� T��������7��� [�����T������� t�����!��W�� {�:�^p� �A�e � $��Z�~/� +/���$/�/p/�/ D/�/h/�/�/�/'?�/ K?�/o?
?�?.?@?R? �?�?�?O�?5O�?YO �?VO�O*O�ONO�OrO �O�O�O�O�OU_@_y_ _�_8_�_\_�_�_�_ o�_?o�_co�_o"o \o�o�o�o|o�o) �o&_�o��B �fx��%��I� �m����,���Ǐb� 돆����3�Ώ��� ,���x���L�՟p��� ����/�ʟS��w��x���ϓ�3 1�� H�Z������6�<�Z� ��~��{���O�ؿs� ���� ϻ�Ϳ߿�z� eϞ�9���]��ρ��� ߷�@���d��ψ�#� 5�G߁�������*� ��N���K����C� ��g��������J� 5�n�	���-���Q��� ������4��X�� Q���q� ��T�x �7�[m�/ />/�b/��/!/�/ �/W/�/{/?�/(?�/ �/�/!?�?m?�?A?�? e?�?�?�?$O�?HO�? lOO�O+O=OOO�O�O �O_�O2_�OV_�OS_ �_'_�_K_�_o_�_�_ �_�_�_Ro=ovoo�o 5o�oYo�o�o�o�o <�o`�oY� ��y��&��#� \�������?�ȏ����4 1�˯u��� ��?�*�c�i���"��� F����|����)�ğ M�����F�����˯ f�﯊�����I�� m����,���P�b�t� �����3�οW��{� �xϱ�L���p��ϔ� ߸������w�bߛ� 6߿�Z���~����� =���a��߅� �2�D� ~��������'���K� ��H������@���d� ����������G2k �*�N��� �1�U� N���n��/ �/Q/�u//�/4/ �/X/j/|/�/??;? �/_?�/�??�?�?T? �?x?O�?%O�?�?�? OOjO�O>O�ObO�O �O�O!_�OE_�Oi__ �_(_:_L_�_�_�_o �_/o�_So�_Po�o$o��oHo�olo�oۏ�5 1����o�o�ol W��o�O�s� ��2��V��z�� '�9�s�ԏ������� ��@�ۏ=�v����5� ��Y��}�����۟<� '�`��������C��� ޯy����&���J�� ��	�C�����ȿc�� ��ϫ��F��j�� ��)ϲ�M�_�qϫ�� ��0���T���x��u� ��I���m��ߑ��� �����t�_��3�� W���{������:��� ^�����/�A�{��� �� ��$��H��E ~�=�a�� ���D/h� '�K���
/� ./�R/��/K/�/ �/�/k/�/�/?�/? N?�/r??�?1?�?U? g?y?�?O�?8O�?\O �?�OO}O�OQO�OuO��O�O"_t6 1�%�O�O_�_�_�_ �O�_|_o�_o;o�_ _o�_�oo�oBoTofo �o�o%�oI�om j�>�b�� �����i�T��� (���L�Տp�ҏ��� /�ʏS��w��$�6� p�џ���������=� ؟:�s����2���V� ߯z�����د9�$�]� �������@���ۿv� ����#Ͼ�G����� @ϡό���`��τ�� ��
�C���g�ߋ�&� ��J�\�nߨ�	���-� ��Q���u��r��F� ��j����������� �q�\���0���T��� x�����7��[�� ,>x��� �!�E�B{ �:�^���� �A/,/e/ /�/$/�/ H/�/�/~/?�/+?�/xO?5_GT7 1�R_ �/?H?�?�?�?�/O �?2O�?/OhOO�O'O �OKO�OoO�O�O�O._ _R_�Ov__�_5_�_ �_k_�_�_o�_<o�_ �_�_5o�o�o�oUo�o yo�o�o8�o\�o ��?Qc�� �"��F��j��g� ��;�ď_�菃���� ��ˏ�f�Q���%��� I�ҟm�ϟ���,�ǟ P��t��!�3�m�ί ��򯍯���:�կ7� p����/���S�ܿw� ����տ6�!�Z���~� Ϣ�=ϟ���s��ϗ�  ߻�D������=ߞ� ����]��߁�
��� @���d��߈�#��G� Y�k�����*���N� ��r��o���C���g� ����������n Y�-�Q�u� �4�X�|b?t48 1�?); u��/;/�_/ �\/�/0/�/T/�/x/ ?�/�/�/�/[?F?? ?�?>?�?b?�?�?�? !O�?EO�?iOOO(O bO�O�O�O�O_�O/_ �O,_e_ _�_$_�_H_ �_l_~_�_�_+ooOo �_soo�o2o�o�oho �o�o�o9�o�o�o 2�~�R�v� ��5��Y��}�� ��<�N�`������� ��C�ޏg��d���8� ��\�埀�	�����ȟ �c�N���"���F�ϯ j�̯���)�įM�� q���0�j�˿��� ��Ϯ�7�ҿ4�m�� ��,ϵ�P���tφϘ� ��3��W���{�ߟ� :ߜ���p��ߔ��� A����� �:���� Z���~�����=���a���� �����M�ASK 1���������XNO�  ���� MO�TE  �R_?CFG �Y�����PL_RAN�GUP���OW_ER ��� ��A��*SYS�TEM*P�V9.�3044 �1/�9/2020 �A � ���R�ESTART_T�   , $�FLAG� $D�SB_SIGNA�L� $UP_�CND4��RS�232r �� $COMME�NT $D�EVICEUSE�4PEEC$PA�RITY4OPB�ITS4FLOW�CONTRO3T�IMEOUe6C�U�M4AUXT���5INTERF{ACsTATU��KCH� t $OL�D_yC_SW �'FREEFR�OMSIZ �A�RGET_DIR� 	$UPD�T_MAP"� T�SK_ENB"E�XP:*#!jFA�UL EV!�R�V_DATA�_  $n E��   	$VAL�U�! 	j&GR�P_   �{!A  2 ��SCR	�� �$ITP_��" $NUMΞ OUP� �#TO�T_AX��#DS}P�&JOGLI�FINE_PCdn�OND�%$�UM�K5 _MIiR1!4PP TN?8�APL"G0_EX�b0<$�!� 814�!P=Gw6BRKH�;&{NC� IS �  �2TYP� �2�"�P+ Ds�#;0BS�OC�&R N�5DU�MMY164�"S�V_CODE_O�P�SFSPD_�OVRD�2^L�DB3ORGTP; LEFF�0<G� �OV5SFTJRUNWC!SFpF5%3oUFRA�JTO��LCHDLY7R�ECOVD'� WaS* �0�E0RO���10_p@  � @��S NVE�RT"OFS�@C� "FWD8A�D4A��1ENABZ6�0T�R3$1_`1FD}O[6MB_CM�!zFPB� BL_M��(!2hRnQ2xCV�"�' } �#PBGiW|8A�Mz3\P��U�B�__�M�P�M� �1�AT�$CA� �PD�2��PHBK+!:&aI�O�4 eIDX+bPPAj?a$iOd�7e�U7a�CDVC_DBG"�a;!&�`��B5�e1�j�S�e3��f�@ATIO� ���AU�c� �S�AB
0Y.#0�D���X!� _�:&S�UBCPU%0S�IN_RS�T, 1�N|�S�T!�1$HW_C1�"]q.`�v��Q$AT! � �_$UNIT�4�p>�pATTRI= �r�0CYCL3NE�CA�bL3FLTR_2_FI9a7�c�,!LP;CHK�_�SCT>3F_ƥwF_�|8��zFS8+�R�rCHAGp�py��R�x�RSD�@`'�1E#&7`_T�X�PRO�`@S�EMOPER_0�3Tf��]p� f��P�DI�AG;%RAILAiC�c4rM� LO�04�A�65�"PS�"�2� -`�e�SPR�`S&.  �W�Ctaf�	�CFUNC�2~�RINS_T.!`(�w��� S_� ��0�P�� 	d��W�ARL0bCBLCUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!��8�3�TID�S��!�� $CE_RIYA !5AFDpPC�~��@��T2 �C�9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@HRgDYOL1	PRG8��H��>1(�ҥMUGLSE =#Sw3��$JJJ6BKGFK�FAN_ALML�V3R�WRNY�HGARD�0+&_P "B��2Q���!�5_�@�:&AU�Rk��TO_SBRvb��� �ƺ�pvc�޳MPINF�@�q�)���'REG'd~0V) 0R<�C�1DAL_ \2sFL�u�2$MԐ (�#S��P� `�gśCMt`NF�qsO!NIP�q5P��IPP� 9a$Y��! �"�!�� �o3EG0P��#@��AR� �c��52�����|5AX�E�'ROB�*REMD�&WR�@�1_=݆�3SY�0ѥ0_�S�i�WRI�@�ƅpST�#��0*@� �q!	���3��� B� �At��3�D�POTO�9� �@ARY�#��0!��d�!1FI�0��$LINK��GkTH�B T_����A��6�"/�XY�Z+"9�7G�OFF��@�.�"���B� l����A3$ ��FI�p���4�4l��$_Jd�"(B�,a������8�"q�������Ck6DUtR��94�TURT�!XZ�N����Xx��P��FL/�@s��l��P��30�"Q +1� K
0M:$�5�3]q7�SuD�Sw#ORQɆ�!�����Q7�
�0O[�ND�=#�!�#�1OVE8��M ���R��R��Q�!P.!P! OAN }q	�R����990�  �brJ9V����Lv�!ER1��	8�!E�@n D�A��p�嘕Ă���v�AX�C�"��`�q� s���0~3� ~F�~e�~�~E�~1��~Ҡ{Ҡ� Ҡ�Ҡ�Ҡ�Ҡ� Ҡ�Ҡ�Ҡ�!)oDEBU}s$x�`��삼!R*�AB��a8A2V`|r 
�"�c���%�Q7� 7�173�7F�7e� 7�7E�����.��LAB����yp��cGRO�p��}��PB_ҁ ��1C���ð�6�1���5���6AND��8p�a3���-G �Q����AH�PH�p2�NTd��Cs@VEL؁�}A��F?�SERVEs@��� $����A!�!�@POR}�KP��b�A�B���	���$�BTRQ�
��CH��@
�G��2	��Eb��_  qlb��Q�ERR��RI�P�@�FQTO	Q�� L�}��YV�ĀG�E%�\���CRE�  �,�A�EP
�RA~�Q 2 d�R�7c��T�@ ��$F ׂ��m����BOC��P � 8[COUNT��ќ��SFZN_wCFG�A 4�p%��rT\zs�a�#`p�Jp c%d�� �� MGp+����`�OGp�eFAq����cX8еk�ioQ��'ѴD�p8�Pz���HE�LA�-b }5��B_BAS\�RSR$�`�2�SH��L�!p1�W!p2DzU3Dz4Dz5Dz6Dz�7Dz8�WqROO0���P�1�NL�� ��AB�C
�"pACK��&IN�PT+�W�Up��	�k��y_PU8�,~�|�OU�CP��%��s�Vl���YTPF?WD_KARKQ-�&:PRE�D�P����QUE$�Ā9 )���~���IU��#s/�p��@�/�SEM1�ǆ1�A�aSTYf�tSO����DI�q���Qc��X��_TM>9�MANRQ �/��END��$KEYSWITCH2��G����HE)�BE�ATMz�PE��L�EJR���0x�UF�F���G�S�DO_H�OM��Oz��pEFPR��SbJі��u�C��O��7P�QOV�_M��}�c�IOC�M���1�BsHK�� D,�&�a`	U2R��M��a�r +��FORC*�WARn���� uOM��  @�$�㰰U��P�1��g���e3��4�1.��S�P�OW�Lz��R%�U�NLO�0T�E�D��  �SNuP��S.b 0N��ADDa`z�$S{IZ*�$VA�0~�UMULTIP�r�P���Az� � $��ƒ����SQc�1CFPv�F'RIFr�PSw����ʔf�NF#�ODBUx�R@w������F��:�IAh�����������S"p�� �  �cRTE���SGL.�T�x�&�C`Gõ3a�/�STM�T��`�P����BW<9 0�SHOWh�q7BANt�TPo���@E�����PV�_Gsb �$PaC�0�PoFBv�-P��SP��A�p����PVD��rbw� �+QA002D .ҝ�6ק�6ױ�6׻��6�54�64�74�8*4�94�A4�B4و� 6ׇ17�}�6�F4�  ��@�����Z����t�U1��1��1��1��U1��1��1��1��U1��1��23�2@�U2M�2Z�2g�2t�U2��2��2��2��U2��2��2��2��2��2��33�����M�3Z�3g�3t�3���3��3��3��3���3��3��3��3���3��43�4@�4�M�4Z�4g�4t�4���4��4��4��4���4��4��4��4���4��53�5@�5�M�5Z�5g�5t�5���5��5��5��5���5��5��5��5���5��63�6@�6�M�6Z�6g�6t�6���6��6��6��6���6��6��6��6���6��73�7@�7�M�7Z�7g�7t�7���7��7��7��7���7��7��7��7���7��hbVPv�U�B �@�09r�
o�V���A x� �0R���  ��BM�@RP�`�4Q_�PR�@[U�AR��D�SMC��E2F_�U��=A ��YSL|�P�@ �  � ֲ>g�������iD��VALU>e�pL��A�HFZAID_L����EHI�JIh�$FILE_ ��D�dc$Ǔ�PXCSA�Q� h�0!PE_BLCKz�.RI�7XD_CPUGY!�GY��Ic�O
TUB���R�  � PaW`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q��TJ��U�Q�T�Q�UH`��T`�T@�T2L��_LIz�  ]�pG_OT�P_EDIU�-b�`7c ?bة�pBQh�~�� �TBC2 �! �%�>��P���a�7aFTτ�d݃T�DC�PA�N`�`M0�0�f�a�gTH��U��d�3�gR�q�9�ERVEЃt݃t�	��a�p�` "�X -$EqLE�NЃRt݃Ep�pRA�v��Y@W_AtS14Eq�D2�wMO?Q�	S���pI�.B�A�y��4Ep�{DE�u��LgACE �CCC�.B��_MA��v��w�TCV�:��wT,�;�Z�P���sѨ~��s�J�A�MD����J���uā
�uQq2ѐ���݁l�s�JK��VK�� ����	���J�����JJ�JJ�AAL�<��<�6��2:�5�cm�N1a�m�(,��DL�p_\�Q�0ApCF
�# `�0GROU�@J�Բ���N�`C^�ȐRE�QUIRrÀEBqUu�Aq��$T�p2"��Bp薋a	��d�$ \?@qhAPPmR��CLB
$H`�N;�CLO}`K�S��e`��u
�aI�% �3�M�`�l��'_MG񱥠C �"Pp����&���BRK���NOLD����RTCMO6a�ޭ��J6`�P>��p��p��pPZ��pc��p6+�7+��<����e&� �lr��������PATH���������qx�����%0A��S�CAub��<���INFDrUC�p�q�C�KUM�Y�psP�� ��A q/ʤ�/�E�/��PAYLOA�J{2L�0R_AN�ap�L�Pz�v�jɆ����R_F2LSHRt��LO{�R����|���ACRL_�q �����b�d�H�@B�$H��"�FLE�X>�$�`J�f' P(��o�o+�p�>�Du( : Qcv�p����fe��po��|F1���-瀢�����]�E ��*�<�N�`�r��� ��4�Q�������A�c� ��ɏۏ���T��2�X:A������ ����)�;�?�H�6��Z�c�u�����.`BJ��) ��`��˟ݟ��`�0ATF�𑢀E�L��(a��J�(v��JE۠CTR���A�TN�1�HA_ND_VBB>�ܯ@�* $��F24���d�CSW>�=s���+� $$M �����0ˡ�ڡ������A�@g����AD)��A���@˪A٫AA� ��`P˪D٫�D�PȰG�P�)S�Tͧ�!ک�!N�DY�P9����#%��Fp ���Ѫ���i����������P3�<�E�N�W��`�i�r���J�e,1 ��ԓ� n�5<m��1ASYMص.@	�ض+A������_`��	���D� &�8�J�\�n�Ju�&���ʧC�I��S�_VI�o�Hm��@V_UANVb�@
S+��J� "RP5"R��&T��3TWV �͢���&��ߪU��a/�7�w��`HR`�ta-��QQ�1�D)I��O�T����PN��. ; *"IAA*���$aG�2C2cJ��$��I��P / �� �ME��� Mb�R4AT�PPT@�@� ��ua���PАl@zh�a�iT�@��� $DUMMY}1E�$PS_D�RF�w�$�fn3�FLA��YP����b}c$GLB_T��Uuu`1�� ��EQa0 X(����ST����SBR��PM21_V��T�$SV_ER��O�_@KscsCLpKrA���O'b�PGL�@E�W��1 4��a+$Y|Z|W�s����AN`�  ��sU�u2 ��N��p�@$GIU{}$�q 1�t�p��3 L���v^B�}$F^BE�vNE+AR��NK�F8����TANCK�  ��JOG��� �4� $JOIN�T�����uMSET.��5  �wE�H�� S����� ��6��  MU��?����LOCK_F�O����PBGLV�HGL�TEST�_XM>���EMP�t����r̀$1U�Гr��22���sB,�3���Ҁ,�1Mq�CE���sM� $K�AR��M�STPD�RA�pj�a�VECX��{�e�IU,�41�{HEԀTOOL�ڠ�V�RE��IS�3����6N�A�AC)H���5��O�}cj�d3���pSI.��  @$RAI�L_BOXE���ppROBO��?�~pqHOWWAR*�x��`�ROLM�b B���S��
�5����O_F� !ppHOTML5�Q�����AP�QGU�C�H��7m�
��R
��O��8m��v�z��!p�sOU��9 	tpp(�14A�̀���PO֡%PIP��N��
�ڑS��,�����CORDEaDҀް̠5�XT���q)���P� O4` �: D pOBP!"Ҁ{�j��cp�j�^@$SYSj�A�DR#�Pu`TCH�� ; ,��E�N�RZ�Aف_�t�״�>��PVWV�APa< � �p��r�UPREV_�RT]1$EDI}T�VSHWR��7v;���q�@D�_`#R�+$H�EADoA�Pl�A�$�KE�q�`CPS�PD��JMP��Ld�U� R��d=r�TO�϶I�S#Ci�NE��$_TIC�K�AMX�AS���HN-q> @pt������_GP֜�[�STYѲ�LAOq���Ҩ�?�5
�Gݵ%$���tu=7pS !$Q ��da�e!`�fP�0ևSQUd� ��b�ATGERCy`|�pS�@ �pCp����d�%Oz`mcO�IZ�d�q�e�aP�RM��a8����PU�QH�_DO=�ְXuS��K�VAXIg�f�1�UR� ��$ #�Е��� _�����ET��Pۂ���5�f�F�7g�A�!�1U�d9�2;]��TSR|Al �о���#��5�� #��#�)#�)i�>' i�N'i�^&{����){�H���2��C����C���WOiO{O�D�qSSC�p B hppD1S(�a�`SP`�ATL �I����~�bADDRES��=B'�SHIF��"��_2CH#��I\&p��TU&pI�� C͢CUST}O��AC�TV��IbDȲ,��0�
�
��U�R`E \�����f�7���tC�#	���F���irt�TXSCR�EEl�F�P��T�INA�s�p��tpb����0G T�� fp,⧱eqBp&uᦲ8u�$#�RRO'0R�`��}�!Ce�pUE��GH ��0���`S�qN��RSM�k�UV�0���V~!�PS_�s�&@C�!�)�'C��Cǂ�z"� 2G�0U�E�4Ibvr�&8�G+MTjPLDQ��Rp��z�BBL_�W��`R`J �f�>2O�qJ2LE�U3"��T4RIGH^3B�RDxt�CKGRĦ`�5TW��7�1WIDTH�H����a�a����UIu�E9Y��QaK d�p���A�J�
�4�BAC�KH��b�5|qX`F�OD�GLABS�?�(X`I�˂$UAR(�9@��0^`H4!� L 8�QR�_k��\B_`R�p͂�����HBO�R`M���w0Uj0�CRۂM�LUM�C��� �ERV�\!I�PN�E�4NV`��GE`=B#���]�t�LP�E��E��Z)Wj'XPz'XԐ&Y5$[6$[7$[8	R���3�<����fԑŁS���M�1USR�tO <��^`U�r�rsFO
�rPRI���m����PTRIP��m�UNDO��P�p��`m�4�l�C�#���� �QWB�P7�G �s�Tf�H�RbOS�agfR��:">c��.qR��s�~�b*��!$�	UQ.qS�o�o�#R�)�>cOFF���pT� �cOp 1�R�t/tS�GU��P.q��JsETw�1�SUB*� f�E/_EXE��V��>c�WO>� U�`�^g��WA'��P�qz!@� V_DB�s��p�2SRT�`
�V0�Q�r��OR��u'RAU��tT�ͷr�q_���W |%��͸OWNA`޴$GSRCE � ��D��<\��MPFIA�p��ESPD����� �C���Gƒ�@+�5��!GX `�`�r޴�n��COP�a$��C`_w������rCT�3�q���qƒp���@� Y"SHADOW�ઓ@�?_UNSCA��@���4M�DGDߑ��E�GAC�,Me�G��Z (0NOX�@�D<�PE�B��VW�S�G���![o � ��VEE#��ڒANG�$��c�薴cڒLIM_X �c��c� ����#`��`� 퐾�VF� ��s�VCCjв�\ՒC{�RAlצ���\RpNFA��Z%�E��Z`G� f^0[�C`DEĒ��� STEQ1���@ �ꁻ@I��`+0���p�`����P_A6��r���K��!]�# 1Ҡ�����\�ȫсCPC�@]�DRIܐ\�͑V#Ѐ����D�TMY_UBY�T���c��F!���bY�븲���P_V��y��LN�BMQ1�$��DEY��EXX�e��MU��X�M� US�!���P_AR����P� ߖG��PACIr�ʐf�ᔀ���c�´c���#�EqB��a.2B���Ч^ ܀GΐP����)�D�R~``�_ �0�@3!�1zr	�e�R�SW��p�00��$S�6�O�Q�1A� XӚ#�E�UE��00���C�HKJ�`�@�p���U� �EA�N�ٖp�pX��MR�CV�!a ��@O*��M�pC�	��s����REF*7
��� �����/��P��@��� @��b��֗�_Y��� ���ۣ��Q$3���8��?��$b �����%���Q��$GROU� �c�����ʠ]��I2^0��U` 0_�I,�o V� ULա`��C&�frAaB�?�NT�� �������A���Q��K�L����õ��A���Qr��T a$c t�`3MD�p8�HU���vSA�CMPE �F  _�R r�p@����XS	���GF/�b#d, �&�@M�P^0۰UF�_C !���z �RO h0"+���@���0C��UREB���RI��
IN�p������d��d��ca�IN"E�H�y��0V�a-�걗�3�W����`���C��i�LO��}�z�@0�!�QNSI��݁���c$&�c$&^.�X_PE-YW+'Z_M�ڒW�Iӑ$�" �+R�'rR;SLre �/�IM
`�RE�C7�Gd�۰�̵ҭ�q��� �u��Ȑ���`���S_P�VnP *��IA�vf �~pHkDR�p�pJO�P���$Z_U�P��a_LOW��5�1J�dA��LINubEP?�tc_i�1�1���@�G1@��V��xg 5X�P�ATHP X�CACH$�]E��yI��A��{�C)�ID3F�A�ETD�H��$H�O�pղb@�{��d6�F�����p�PA3GE�䁀VP�°��(R_SIZ��2TZ�3�-X�0U�q�MP\RZ��IMG���sAD�Y�MRE���R7WGP��8�p��ASYNBUF�VRTD�U�T7Q�LE_2D-��U�J�`CҡU1��Qu���UECCU��VE�M��]EDb�GVIR�C�Q�U�S�B�Q�L�A��p�NFOUN^_�DIAG�YRE�GXYZ�cE�W� �h8�dpqa`T��2IM�a�V|be��EG/RABB��Y�aЗLERj�C4���FC-A�6504x��7u��� BE��h'�>`�CKLAS_@l�8BA��N@i  G��IT��� @ݲմ$BAƠwj �!q�eb��uTYSp�H����2B��I�t:b�f��B)�gEVE����PK��؂fx��GI�pNOt��2�\r_HO��>��k � ���
8�Pi�S�0ޗ���RO�ACCEL�?0=���VR_�U�7@�`��2�p��ARF��PA��̎K�D���REM_But M�rJMX �l�t>�$SSC�Uk� #���QN@m �� �S�P�NS����VLEX�vn =T�ENAB 2¼W@��FLDRߨF�I�P�t�ߨ(Ğ���2P2HFo� ���V
Q MV_PI��8T@�H���F@�Z� +�#��8�8#��sGAB���LOO󣎔�JCBx��w"SC�ON(P�PLANۀ�Dp�3F�d�v�9PէM��Q ;����SM0E�ɥ�8ɥWb 72$`<�8T��,`�RKh"ǁVANC���@AR_Ou N@p (�-#<#c��c�2 w�A/�N@q 4������`	�^�� w�N@r hn���1�^�&OFF`|�p��`��`�DEA�
��P,`SK�DMP6V{IE��2q w���@���rs < {���4���r{7���D��Ȭ!CUS�T�U��t $�G�TIT1$sPR\��OPTap� ��VSF�йsuB�p�0`r&��1SMOwvI�|�ĄYJ�����eQ_WB��wI���� @O3��@�XVRxx�mr��T��
�Z�ABC��y �op����)�
}qZD�$�CSCH��z Lu����`�2�%PC ��7PGN ��<�<�A��_FUNH��@�)P�ZIPw{,I��LV,SL��~�}��ZMPCF���|��E����X�DMY_LNH�=�C�� ~��} $�A�� ]�CMCM� C�,SC&!��P�� �$J���D Q�������������a_�Q,2����UX�a>\�UXEUL��a ������(�:�(�J���FTFL��w�7�Z�~Zp+�T6����Y@Dp�  8 $�R�PU��> EIGH����?(�iֱ�q�0��et� �a�����$B�0�0@�}	�_SHIFD3�-�RVV`Fcв�		$5��C�0��&!������b
�sx�uMD�TR��V̱���SPH���!�� ,������� ��4A�RYP��%������%��"��%!  �H�(UN0���"�2 �����ɐ�q0�GSPDak����P��O�����0��첱��"!NGVER`q �iw+I�_AIRPURG�E  i  �i/�F`E�Tb� ��+  � h2I�SOLC  �,"�"�!!�%�²P+�_/*OB��D�m�?@�!�H771   34n?�?�9� `�E/#z�)x� S232��� 1i� L�TEk@ PENDA�341 1D�3<*? �Mainten�ance Con%s B�? F"O,DNo UseM JOOnO�O�O�O�O2��2NPO;� 1�9%�1CH=� 9�-Q		9Q_?!UD1:___�RSMAVAIL�/�/%�A!SR  �+��H�_�P�1�TVAL.&����P(.�YVL�}� �2i�� D��P 	�/_oUQ No�orci�o�g�o�o �o�o�o*,> tb������ ���:�(�^�L��� p�������܏ʏ �� $��H�6�X�~�l��� ��Ɵ���؟����� D�2�h�V���z����� ���ԯ
���.��R� @�b�d�v�����п�� �����(�N�<�r��i�$SAF_D?O_PULS. j0Qp����CA� ��/%�&0SCR ��` �X�
�0�0
	14�1IAIE���b vo$�6� H�Z�l�~�ߢߴ��߰�������HS"��2%�����d1�(��8�rb��� @��"k�}���T�h� �J`���_ @��T7 �����#�~0�T D��0� Y�k�}����������� ����1CUg�y�O�Ef�p����  �5�;�o�� 1p��U�
�t���Di�������
  � ��*������ gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O7O<A���`OrO�O�O �O�O�O�O�O?O�_ ._@_R_d_v_�_�_�_�_�Q _�R0MJ To!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏJO��'�9�K� ]�o�������_ɟ۟ ����#�5�G�Y��_ �U�_�ҙ�����ϯ� ���)�;�M�_�m� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�;�?� q߮����������� ,�>�P�b�t�������������������Y��	�1234567�81h!B�!����F��� ��������������  ��;M_q ������� %7I[l*� ������// 1/C/U/g/y/�/�/�/ n��/�/	??-??? Q?c?u?�?�?�?�?�? �?�?O�/)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_O_ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �op_�o�o�o/ ASew���� �����o+�=�O� a�s���������͏ߏ ���'�9�K�]�� ��������ɟ۟��� �#�5�G�Y�k�}����������s�կ��w���0�L�CH�  Bpw�   ��=�2�� �} =�
~���  	�o�@ί��ǿٿ���r������@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖ�%� ����������&�8� J�\�n��������������"�Q�*�(����;�<M���D�~��  �]��w�*�Z򛱛�t C d�����*�`*���$SCR_GR�P 1 *P� 3� � }�*� 6��	 �
��<�+�*�'UC|@�Y�y�yD� W��!�y�	M-�10iA/7L �12345678k90��� 8���MT� � �
��	L��	Č� N
���Y���Dy�
M_	P������ ,���H�
 � ��1/@A/g/y/H���!T/�/P/�/3��+\���/B�S��,?�*2C4&Ad�R?  a@s�j5N?�7?��7�&2R��?}:&F@ F�`�2�?�/�? �?OO-OSO>OwObO �O=j1�2�O�O�O�O�DB��O�O;_&___ J_�_n_�_�_�_�_�_ o�_%o�5j�eSgxo6���uo�o�b�1�B�|3�oh0�4j96j9B� w�$0Y̯@HtA�Nhcu$�/�%pp�drsqA ����z�q�x�� �� (&� *�2�D�V�oz�e��������ECLVL ; ����iqp�Q@��L_DEF�AULT ���s�փH�OTSTR�qq���MIPOWER�F��H���WF�DO� �RVENT 1Ɂ�Ɂ� L!D?UM_EIP������j!AF_I�NE‧���!FIT}�֞����!-/�� ��F�!�RPC_MAIN�G�)��5���Y�VI�Sb�t����ޯ!�TPѠPUկ��d�ͯ*�!
PMON?_PROXY+���Ae�v��D���fe��¿!RDM_S�RVÿ��g���!#R,*ϑ�h��Z�K!
[�M����iI����!RLSYN�C����8����!�ROS|���4���>�!
CE�MOTCOM?ߓ�k-����!	S�CONSd�ߒ�ly���!SҟWASRCݿ��m���"�!S�USB�#n�n�!S#TMC��o]�� ���ѳ����,����P�V�ICE_KL� ?%d� (%�SVCPRG1S�����2�������oD����4������5D��6;@��7c h�����9����%������� ��0����X��� ��-���U���} ��� /���H/�� �p/���/��F�/ ��n�/��?�� 8?���`?��/�?�� 6/�?��^/�?��/X� j��q���#OhO��lO �O{O�O�O�O�O�O�O  _2__V_A_z_e_�_ �_�_�_�_�_�_oo @o+odoOo�o�o�o�o �o�o�o�o*< `K�o���� ���&��J�5�n� Y���}���ȏ���^�_DEV d���MC:�4����GRP �2d�
@�bx� 	� 
 ,V�ȡ�s�Z����� �������ߟ�� @�'�9�v�]�������@Я����۫Y��
@�ܯI�1�4�]��� j�����˿F�Ŀ�� %�7��[�B��f�x� ���!���A����ۿ D�+�h�Oߌ�s߅��� ������
���@�'�d�v��	y��^��� ��������%��I�0� Y��f�����8����� ������3��T7]�e�����)� �
�.@�dK �o��!�9���!/G/���R/ �/�/�/�/�/"�/�/ ??C?*?<?y?`?�? ��?�?�?�?�?�?-O OQO8OaO�OnO�O�O �O�O�O_�O)_;_"_ __�?�_�_L_�_�_�_ �_�_o�_7oo0omo To�oxo�o�o�o�o�o !x_E�oU{b �������� /��S�:�w�^�p������я�d �XƿZI6 r���@Z��0�+�A����d�BjBA�=��������B����AZ.�A����+�A.��Q�B�����5\��i6�A��u��'��ǎ%�Ꮛ�%�PEGA_BAR�RA_ESTEI�RA����X�T����?=��=�X��7
�?��>�A����?������&����������AxP��f���U�'A�j���´�B��:�<�3�����jB]+a��T��%�T�腯d�ʐ���>�p�c?��7�Գ�T@6��A�_���0n�����·�Ak���۸I�K9�FA�G�����B!v,�-���C3�����pBM�>�#�b��(�Y�������HX��?L!���Q��B���AJߤ�Xk�@f�D3��O�A���������Yw���.B��B�;��C�H�z�B�?���6���-Ϙ������n��=]����V@����?,����Ö� վ���eAk�������OY�A��ㇾ��AB��J�;%�C$�4�aƿBXZ�9���
���ߘ��~��� �ԭ(��?^_��-\¯ԡ���گ���+������������ߔ�mᢧ��*נ�6�C>�ԯb���z���
��BM����s��x�U<~�߯7@6|=��C��$�6��� N�@���b�G���L��}������x7���~K@����V�+A>r�rF���������Y@+�@��<B��|�A��F����B)���,o�?ɇ���~0��0~�6�Z� Q������������Aߍ�]ܖ�A����ܺ����2[�����>�ȥA���=�³�NB ��$�w?�d�j��to�7\��
�.�%��Z�����A������*�@Ve��B� ������YN�#���BD�	����9A����gB#
q��3��C4#���,?[BVM����COLO�CA_PRENS�����&//J/ 8/n/\/~/�/�/ �/�/�/ ??D?2?T? �/�/�?�/z?�?�?�? �?O
O@O�?gO�?0O �O,O�O�O�O�O�O_ ZO?_~O_r_`_�_�_ �_�_�_�_2_oV_�_ Jo8ono\o�o�o�o�o 
o�o.o�o"F4 jX��o��~� z���B�0�f�� ���V�����Џҏ� ��>���e���.��� ������̟Ο���X� =�|��p�^������� ��ȯ�D��T��H� 6�l�Z���~�����ۿ ���Ϡ��D�2�h� Vό�ο���|����� 
����@�.�dߦϋ� ��T߾߬�������� �<�~�c��,��� ��������D�)�;� �����\��������� ���@���4"D FX�|���� ��0@BT ����z��/ �,//</���/� b/�/�/�/�/?�/(? j/O?�/?�??�?�? �?�?�? OB?'Of?�? ZOHO~OlO�O�O�O�O O�O>O�O2_ _V_D_ z_h_�_�_�O�__�_ 
o�_.ooRo@ovo�_ �o�ofo�obo�o�o *N�ou�o>� ������&�h M�����n������� ��ȏ��@�%�d��X� F�|�j��������,� ��<�֟0��T�B�x� f���ޟï������� �,��P�>�t����� گd�ο�����(� �Lώ�sϲ�<Ϧϔ� �ϸ�������$�f�K� ���~�lߢߐ��ߴ� ��,��#�������D� z�h��������(� ���
�,�.�@�v�d� ������ ������� (*<r����� b����$ z�q�J��� ���/R7/v / j/�z/�/�/�/�/�/ */?N/�/B?0?f?T? v?�?�?�??�?&?�? OO>O,ObOPOrO�O �?�O�?�O�O�O__ :_(_^_�O�_�_N_p_ J_�_�_�_o o6ox_ ]o�_&o�o~o�o�o�o �o�oPo5to�oh V�z����( �L�@�.�d�R��� v������$���� �<�*�`�N���Ə�� �t�ޟp����8� &�\�����L����� گȯ����4�v�[� ��$���|�����ֿĿ ��N�3�r���f�T� ��xϮϜ������� ���Ͼ�,�b�P߆�t� ������ߚ����� �(�^�L���ߩ��� r����� �����$� Z������J������� ������b���Y�� 2�z����� :^�R�b� v����6� *//N/</^/�/r/�/ ��//�/?�/&?? J?8?Z?�?�/�?�/p? �?�?�?�?"OOFO�? mOO6OXO2O�O�O�O �O�O_`OE_�O_x_ f_�_�_�_�_�_�_8_ o\_�_Po>otobo�o �o�o�oo�o4o�o( L:p^��o�o �� ��$��H� 6�l�����\�ƏX� ֏��� ��D���k� ��4�������ҟ�� ��^�C����v�d� ��������ί��6�� Z��N�<�r�`����� �����󿪿̿��� J�8�n�\ϒ�Կ���� �����������F�4� j߬ϑ���Z��߲��� �������B��i�� 2������������ J�p�A����t�b��� ��������"�F��� :��Jp^��� ���� 6$ FlZ����� ��/�2/ /B/h/ ��/�X/�/�/�/�/ 
?�/.?p/U?g??@? ?�?�?�?�?�?OH? -Ol?�?`ONOpOrO�O �O�O�O O_DO�O8_ &_\_J_l_n_�_�_�O �__�_o�_4o"oXo Foho�_�_�o�_�o�o �o�o0T�o{ �oD�@���� �,�nS�����t� ��������Ώ�F�+� j��^�L���p����� ��ܟ��B�̟6�$� Z�H�~�l����ɯۯ ��������2� �V�D��z��������$�SERV_MAI�L  �����ʴOUTPUT�ո�@�ʴRV 2j� � � (r�������=�ʴSAV�E���TOP10� 2� d 6 rƱ���� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t������n�YPY��F�ZN_CFG f��=���J���GRP 2���g� ,B  � A �D;� �B �  B4~=�RB21I�oHELL��f�e�)�*�=�����%RSR��� ���&J5 G�k�������.�  ���/>/P/"\/ b�X/z"{ �U'
&"2�dh,g-�"E�HK 1S �/�/�/�/#?L?G? Y?k?�?�?�?�?�?�?��?�?$OO1OCO?OMM S�OD�FTOV_ENB�մ�e��"OW_R�EG_UI�O�IMIOFWDL~@��N�BWAIT��B�)��V��F��YTIM�E���G_VA԰_�A_�UNIT�C~Ve�L]C�@TRY�Ge��ʰMON_AL�IAS ?e�I%�he��oo&o8o Fj�_io{o�o�oJo�o �o�o�o�o/AS ew"����� ���+�=��N�s� ������T�͏ߏ�� ���9�K�]�o���,� ����ɟ۟ퟘ��#� 5�G��k�}������� ^�ׯ�����ʯC� U�g�y���6�����ӿ 忐����-�?�Q��� uχϙϫϽ�h����� ��)���M�_�q߃� ��@߹������ߚ�� %�7�I�[����� ����r������!�3� ��W�i�{���8����� ��������/AS e�����| �+=�as ��B����/ �'/9/K/]/o//�/ �/�/�/�/�/�/?#? 5?�/F?k?}?�?�?L? �?�?�?�?O�?1OCO UOgOyO$O�O�O�O�O �O�O	__-_?_�Oc_ u_�_�_�_V_�_�_�_�ooc�$SMO�N_DEFPRO�G &����Aa &�*SYSTEM*�obg $JO�0dRECALL �?}Ai ( ��}>copy m�d:pickup�_barra_e�steira.t�p virt:\�temp\=>1�0.109.3.�23:211520bo�o�o	w}<�o�`torno�o�n�o�k}y5vlace1C�bS����};usumir +��i�k�}��v>�cprens�oG�Z������7|��Ï��bՏf�x���=�furad��<��o������v%�sem_recep1���ʟ`Z�l�~����fco-��?�Q����� }:�udrop*�defeit5�ɯدi�d{��8�.�_15��ɏW��������_2���ſ׿h�z���_33�E�W������p�frs:orde�rfil.dat~��mpback�ϠV���i�{��.tb:*.*2���M�������t2x�:\ ��'��S���f�x��3�a%�7�N�R������� }
xyz�rate 61 ������]�o�������=�6:15300 ;�M�����t�tpdisc 0��0 ����\n���tpconn 0 &8J� ���$߭߮��f x�ߝ�8��L�� /��9����a/s/ �/��)/;/��Q/�/�/ ?p�o�o��K\?n? �?�%9?��?�?�? ���?���?dOvO�O ��?9O�ZO�O�O�? �����OXOi_{_ � 7_?/V_�_�_����/_ �_U?eowo
o���Ao So�o�o�����o�o as��*�?�Y ���ϡ����h� z���1�C�U���� ��������ӏd�v��� -��DX����������֟g�y�����$SNPX_AS�G 2������� ��S%���Я  ?����PARAM ����� ��	��PӤ0�Ө$������O�FT_KB_CF�G  ӣ����O�PIN_SIM + ���}����������RVNOR�DY_DO  �)�U���QSTP/_DSBi��Ͼ��SR ��� � &#�D�O��O�:�TOP_ON�_ERRʿ��o�P_TN ������A��RIN�G_PRMy�ܲV�CNT_GP 2���!���x 	 ����0��#��Gߔ��VD��RP 1��"�8Ѩ�*߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�}�z����������� ����
C@Rd v������	 *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? [?X?j?|?�?�?�?�? �?�?�?!OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLosopo�o�o �o�o�o�o�o 9 6HZl~��� ����� �2�D��V�`�PRG_CO7UNTJ���{�'ENB��}�M��L����_UPD 1>'�T  
k��� ���"�K�F�X�j��� ������۟֟���#� �0�B�k�f�x����� ����ү������C� >�P�b���������ӿ ο����(�:�c� ^�pςϫϦϸ����� �� ��;�6�H�Z߃� ~ߐߢ���������� � �2�[�V�h�z�� �����������
�3� .�@�R�{�v������� ������*S�N`r���t�_INFO 1��Ҁ� 	 ���3���)X@�>���L9 C w��Bb?	�;ӛ�8����,,M�A�@�>>�`� AoB @{w� ?�� >�@���a ����C�Tp���1VC3����"��3������YSDEBU�G��퀍dՉ�S�P_PASS���B?+LOG u���  � 9a�  �с�UD1:\;$<�<"_MPCA-�H�/�/�x!�/ �~�&SAV D)`��%d!|"�%�(�SV�+TEM_T�IME 1D'��� 0   ����
�',5M7MEMBK  셂сd d/�?�?�<wX|Ҁ� @�?C�O:OJLOmORzI�J�%@p1 �O�O�O�O"3 __$_06_H_Z_l_ �n_�_ �_�_�_�_�_�_o"o\�e1oVohozo�o�o �o�o�o�o�o
. @Rdv���O5SK�0�8���?����F+� ��H2�OJ�AJ� ��`��A\O����(�O"�Oяb�ݏ���p�O�  ` 	� ��0p�Z�l�~� r_���9�Ο������$�C�7og�y� ��������ӯ���	� �-�?�Q�c�u�����������T1SVG�UNSPD%% '�%��2MOD�E_LIM �a9"ܴ2�	� �D-۵ASK_OP�TION �9!�F�_DI ENB�  �5%f�BC�2_GRP 2!��u#o2��XB��C����ԼBCCFG 3#��*< #6���U�?H�3�E�~� iߢߍ��߱������  ��D�/�h�S��w� ��������
���.�@�R�=�v�����t� ��u�����c���	 B-f�.��4[ � ������  02Dzh��� ����/
/@/./ d/R/�/v/�/�/�/�/ �(���/?&?8?J?�/ n?\?~?�?�?�?�?�? �?O�?4O"OXOFOhO jO|O�O�O�O�O�O�O __._T_B_x_f_�_ �_�_�_�_�_�_oo >o�/Voho�o�o�o(o �o�o�o�o(:L p^����� ��� �6�$�Z�H� ~�l�������؏Ə�� � ��0�2�D�z�h� ��To��ȟ���
��� .��>�d�R������� z�Я�������(� *�<�r�`��������� ޿̿���8�&�\� Jπ�nϐϒϤ����� �ϴ��(�F�X�j��� ��|ߞ��߲������ ��0��T�B�x�f�� ������������� >�,�N�t�b������� ����������:( ^�v����H ���$HZl :�~����� ��2/ /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?P?R?d?�?�? �?t�?�?OO*O�? NO<O^O�OrO�O�O�O �O�O�O__8_&_H_ J_\_�_�_�_�_�_�_ �_�_o4o"oXoFo|o jo�o�o�o�o�o�o�o �?6Hfx� �������v&���$TBCSG_�GRP 2$�u��  ��&� 
 ?�  Q�c�M���q���������ˏ��*�1�&~8�d, �F��?&�	 HCA������b��CS�B�I������V�>��ͪ�n��쌟ԝB��333,��Blt�����r�AÐ�fff:�L�.�C����l�?����G�w�R���A&��̧�����@��I��-���
�X��u�@�R�����̻������	V3.00>I�	mt7����*� �%��ֶY�_�@ff&� &��H�� N� �O� ; ����� ϏϬ��*�J21�'8���Ϥ�CFG )��uB� E�������d���#��#�I�W��pW�}� hߡߌ��߰������ ��
�C�.�g�R��v� ��������	���-� �Q�<�u�`�r����� ������I�cp" 4��gRw��� ���	-?� cN�r��&�� ����/</*/`/ N/�/r/�/�/�/�/�/ ?�/&??J?8?Z?\? n?�?�?�?�?�?�?O �? OFO4OjOXO�O�O `�O�OtO�O_�O0_ _T_B_x_f_�_�_�_ �_�_�_�_�_,ooPo boto�o@o�o�o�o�o �o�o�o(L:p ^������� � �6�$�F�H�Z��� ~�����؏Ə���� 2��OJ�\�n������ ��������
�@� R�d�v�4��������� ί����ү(�N�<� r�`���������ʿ̿ ޿��8�&�\�Jπ� nϐ϶Ϥ��������� "��2�4�F�|�jߠ� �����߀��� �߼� B�0�f�T��x��� ����������>�,� b�P���������v��� ����:(^L �p�����  �$H6lZ| ������/� / /2/h/�߀/�/�/ N/�/�/�/
?�/.?? R?@?v?�?�?�?j?�? �?�?�?O*O<ONOO O�OrO�O�O�O�O�O �O _&__J_8_n_\_ �_�_�_�_�_�_�_o �_4o"oXoFoho�o|o �o�o�o�o�o�/$ 6�/�oxf��� �����,�>�� �t�b�������Ώ�� 򏬏��&�(�:�p� ^���������ܟʟ� � �6�$�Z�H�~�l� ������دƯ��� � �D�2�T�z�h��� Jȿڿ������
�@� .�d�Rψ�vϬϾ��� �Ϡ������*�`� r߄ߖ�Pߺߨ����� �����&�\�J�� n������������ "��F�4�j�X�z�|� ������������0 B�Zl~(�� �����,P bt�D�������   #� &0/"�$T�BJOP_GRP� 2*��  ?�&i	H"O#,V,��w�� �� �=k%  Ȫ �� �� �$ �@ g"	 �CA���&��SC���_%g!�"G���"k��/�+=��CS�?ϙ�?�&0%0CR  B4�'??J7�/^�/?333�2Y&0<}?�:;��v 2�1)�0-1*20�6?�?�20��7C�  D��!�,� BL���OK:�Z�Bl�  @pB@�� s�33C�1 �?gO ' A�zG�2jG�&�)A)E�O�J;��>|A?�ff@U@�1�C�Z0zjO�Oz@����U�O�$fffx0R)_;^;xCsQ?ٶ4)@�O�_tF�X�_J\EU�_�V:�t	-�Q(B�*@�Ooh �&-h$oZGLo6oDoro �o~o8o�o�o�o�o 3�oRlVd���V4�&`�q�%	�V3.00m#'mt7A@�s*�l$�!�'� E���qE���E��]\E�HF�P=F�{F*�HfF@D�FW��3Fp?F��MF���F��MF��F��şF��F��=F���G��G.8�C�W�RD3l)D���E"��E�x�
E��E��,)FdRF�BFHFn� F���F��MF��ɽF�,
G�lGg!G�)�G=��G�S5�GiĈ;��
;�o�|U& : @Xz&/T��&"�?�0��&=;-ESTPARS  (a E#�HRw�ABLE ;1-V) @�#�R�7� � �R�BR�R�'#!R�	R�E
R�R���!R��R�R���RD	I��`!��ԟ���
�r�Oz����������̯ޮ��Sx�^#  <�����ÿտ���� �/�A�S�e�wωϛ� �Ͽ�������;-w�{� _"��6��1�C�U����%�7�I�[����N�UM  �*`!� $  ��m����_CFG .����!@H IMEBF_TT}���^#��G�VE10m�H�]�G�R 1/��' 8�" �� �A�  ����� ������� �2�D�V� h�z������������� /
e@Rhv ������� *<N`r�� ����'///]/ 8/J/`/n/�/�/�/�/�r���_��t�@~��t�MI_CHAN�S� ~� !3DBGLVLS�~�s�$0�ETHERAD �?��w0�"���/�/�?�?l�$0RO�UTq�!�!��4�?�<SNMAS�Kl8~�}1255.2E�s0OBOTO�st��OOLOFS_D�I}��%V9ORQCTRL 0���#��MT�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo&l�O�Io8omoq�PE_D�ETAIJ8�JPG�L_CONFIG� 6�ᄀ�/cell/$C�ID$/grp1�qo�o�o/壀 �?Zl~���C ���� �2��V� h�z�������?�Q�� ��
��.�@�Ϗd�v� ��������M����� �*�<�˟ݟr���������̯@�}a��� &�8�J�\���^o��c��`���˿ݿ��� Z�7�I�[�m�ϑ� � �����������!߰� E�W�i�{ߍߟ�.��� ���������A�S� e�w����<����� ����+���O�a�s� ������8������� '9��]o�� ��F���# 5�Yk}������`�User View �i�}}1234567890�//,/�>/P/X$� �cx/���2�U�/�/�/�/ ??s/�/�3�/b? t?�?�?�?�??�?�.4Q?O(O:OLO^OpO�?�O�.5O�O�O�O@ __$_�OE_�.6�O ~_�_�_�_�_�_7_�_�.7m_2oDoVohozo�o�_�o�.8!o�o�o�
.@�oagr �lCamera��o����� �ޢE�*�<� N��h�z��������I  �v�)��$� 6�H�Z�l�������� ��؟���� �2�Y��vP9ɟ~������� Ưد���� �k�D� V�h�z�����E�W�I 5����� �2�D�� h�zό�׿�������� ��
߱�W�ދ��X�j� |ߎߠ߲�Y������� E��0�B�T�f�x�� �ulY���������
� ���@�R�d������ ����������W� iy� .@Rdv�/�� ���*< N��W��i���� ����/*/</� `/r/�/�/�/�/as9F/�/??1?C?U? �f?�?�?D/�?�?�?��?	OO-O�j	�u0 �?hOzO�O�O�O�Oi? �O�O
_�?._@_R_d_ v_�_/OAO�p�{,_�_ �_oo)o;o�O_oqo �o�_�o�o�o�o�o �_�u���oM_q� ��No���:� %�7�I�[�m�NEa� ���ˏݏ���� 7�I�[���������� ǟٟ����ͻp�%�7� I�[�m��&�����ǯ �����!�3�E�� ��9�ܯ������ǿٿ 뿒��!�3�~�W�i� {ύϟϱ�X�����H� ���!�3�E�W���{� �ߟ������������<���  ��L� ^�p���������x�� ��   "� *�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/��  
��(  ��@�( 	  �/�/�/�/�/? ?6? $?F?H?Z?�?~?�?�?t�?�*2� �l� O/OAO��eOwO�O�O �O�O��O�O�O_TO 1_C_U_g_y_�_�O�_ �_�__�_	oo-o?o Qo�_uo�o�o�_�o�o �o�o^opoM_ q�o������ 6�%�7�~[�m�� �������ُ���D� !�3�E�W�i�{�ԏ ��ß՟�����/� A�S���w�����⟿� ѯ�����`�=�O� a�����������Ϳ߿ &�8��'�9π�]�o� �ϓϥϷ��������� F�#�5�G�Y�k�}��� �߳���������� 1�C�ߜ�y����� ��������	��b�?� Q�c������������ ��(�)p�M_�q������0@ A�������� ��#frh:�\tpgl\ro�bots\m10�ia4_7l.xml�Xj|��������.�� /1/C/U/g/y/�/�/ �/�/�/�/�//?-? ??Q?c?u?�?�?�?�? �?�?�?
?O)O;OMO _OqO�O�O�O�O�O�O �OO _%_7_I_[_m_ _�_�_�_�_�_�__ �_!o3oEoWoio{o�o �o�o�o�o�o�_�o /ASew��� ����o��+�=� O�a�s���������͏�ߏ�I |�<<  ?��4��,�N� |�b�������ʟ�Ο ���0��8�f�L�~�@��������������(�$TPGL_�OUTPUT �9����� $�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}ϏϡϠ������$����2�345678901��� �2�D�V�^� ���υߗߩ߻����� w����'�9�K�]���}g��������o� ����1�C�U�g��� u�����������}��� -?Qc��� ������) ;M_q	�� �����%/7/I/ [/m///�/�/�/�/ �/�/�/?3?E?W?i? {??%?�?�?�?�?�? O�?OAOSOeOwO�O !O�O�O�O�O�O_�O~� $$Ӣ ��OW=_o_a_�_�_�_ �_�_�_�_�_#ooGo 9oko]o�o�o�o�o�o �o�o�oC5g}���������}@��"�� ( 	 iW�E� {�i�����Ï��ӏՏ ���A�/�e�S��� w��������џ��� +��;�=�O���s�����Ƹ  <<\ޯ�)�ͯ�)� �M�_���ʯ����<� ��ؿ��Ŀ� �~�$� V��BόϞ�x����� 2ϼ�
ߤ���@�R�,� v߈���p߾���j��� ����<�߬�r�� ��������`� &�8���$�n�H�Z��� �����������"4 Xj��R��L ����|T f ��v��0 B//�&/P/*/</ �/�/��/�/h/�/? ?�/:?L?�/4?�?? n?�?�?�?�? O^?�? 6OHO�?lO~OXO�O�O O$O�O�O�O_2__ _h_z_�O�_�_J_�_��_�_�_o.o��)�WGL1.XML��cm�$TPOF?F_LIM Š�p����qfNw_SVy`  �t��jP_MON �:���d�p��p2miSTRTC�HK ;���f�~tbVTCOMP�AT�h*q�fVWV_AR <�mMx.�d  e�p��bua_DEFPROG %�i�%COLOC�A_MESA_IRVISI�`�r?ISPLAY�`�n��rINST_MSwK  �| �z?INUSER �t�LCK)��{QUI�CKME�pO��rS7CREl���+r?tpsc�t)�Ї����b��_��ST�z�iRACE_C_FG =�iMtu�`	nt
?��?HNL 2>�z���T{ zr@�R�d�v����������К�IT�EM 2?,� ��%$12345�67890�%� � =<�C�U�]� G !c�k�wp'� ��ns�ѯ5����k� �����j�ů��鯕� ��A�1�C�U�o�y�� ��I�oρ�忥�	�� -ϧ�Q���#�5ߙ�A� ������e߳������ M���q߃�L��g��� �����%�w� �[� ��+�Q�c���o��� �����3���{� ;������G_��� �/�Se.�I �m��� =�a/3/��� ���k//�/�/�/ ]/?�/�/�/?�/u? �?�??�?5?G?Y?�? +O�?OOaO�?mO�?�? �OO�OCO__yO+_ �O�Ox_�O�_�O�_�_ �_?_�_c_u_�_o�_ Wo}o�o�_�oo)o;o �o�oqo1C�oO�o �o��%��[���Z��S�@|��_��  ے�_� ����y
 �Ï�Џ���UoD1:\���q��R_GRP 1A� �� 	 @�pe�w�a���������ߟ͞����ّ��>�)�b�M�?�  }���y�����ӯ�� ����	��Q�?�u��c���������Ϳ�	�-���o�SCBw 2B{� h� e�wωϛϭϿ��������e�UTORIAL C{��@�j��V_CONFIG D{����������O�OUTPUT �E{����� ������%�7�I�[� m���������� ����%�7�I�[�m� ��������������� !3EWi{� ������� /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ ��/??'?9?K?]? o?�?�?�?�?�?�/�? �?O#O5OGOYOkO}O �O�O�O�O�O�?�O_ _1_C_U_g_y_�_�_ �_�_�_�O�_	oo-o ?oQocouo�o�o�o�o �o�_�o);M _q������ yߋ����-�?�Q�c� u���������Ϗ�� �o�)�;�M�_�q��� ������˟ݟ� �� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ���
��/�A�S� e�wωϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ���������1C Ugy����� ��	-?Qc u�������|/�x���$/ 6/ !/a/��/�/�/ �/�/�/�/??'?9? K?]?�?�?�?�?�? �?�?�?O#O5OGOYO kO|?�O�O�O�O�O�O �O__1_C_U_g_xO �_�_�_�_�_�_�_	o o-o?oQocot_�o�o �o�o�o�o�o) ;M_q�o��� �����%�7�I� [�m�~������Ǐُ ����!�3�E�W�i� z�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9��K�]�o�~��$TX�_SCREEN �1F8%  �}�~���������
����m&��\� n߀ߒߤ߶�-�?��� ���"�4�F��j��� ����������_�� ��0�B�T�f�x���� ����������� >��bt���� 3�W(:L ^������� �e/�6/H/Z/l/�~/�//�/�$UA�LRM_MSG k?����� �/ ���/�/)??M?@?q? d?v?�?�?�?�?�?�?�O�%SEV  ��-EF�"ECFoG H�����  ��@�  }AuA   Bȁ�
 O���ŨO�O �O�O�O__&_8_J_�\_jWQAGRP 2�I[K 0��	 ��O�_� I_BB�L_NOTE �J[JT��#l������g@�R�DEFPRO� %��+ (%CO�LOCA_MES�A_IRVISION�_%OVoAozo eo�o�o�o�o�o�o�o�@�[FKEYDATA 1K�ɞ�Pp jG����_������z,�(����(POINT M'�(�v@�CROS�}�d�RE�L  T��� C?HOICE]��)��TOUCHUP ׏؏�'��K�2�o� ��h�����ɟ۟����#�5��Y��y���/frh/gu�i/whitehome.pngd�`����Ưدꯀ{�point���0��B�T�f���   �gmacro������ȿڿ�{�gkarel��(�:�L�^�p���clos��ϯϠ����������{�t?ouchup�0ߠB�T�f�x���{�arwrg������� ���߁��)�;�M�_� q����������� ���%�7�I�[�m�� ������������� ��3EWi{� ������/ ASew��r�� ����/!/(E/ W/i/{/�/�/./�/�/ �/�/??�//?S?e? w?�?�?�?<?�?�?�? OO+O�?OOaOsO�O �O�O8O�O�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o �_Goko}o�o�o�o�o To�o�o1C�o gy����P� �	��-�?�Q��u�@��������Ϗj�܋�u�܏�(�s��Q�c�r�,I���A�OINT  ]��~�� OOK Tß��}�NDIREC�ܟ�  CHOI�CE�����UCHUPG�H�s���~��� ��߯�د���9�K� 2�o�V�������ɿ���whitehom����%�7�I�X���poin�ߍϟ�������d�i/look}��(�:�L��^�i�indirec|Ϙߪ߼�����g�choic���� ��2�D�V�h�k�touchup�ߠ���������g�arwrg ��"�4�F�X�j�a��� ����������w� 0BTfx�� �����,> Pbt���� ��/�(/:/L/^/ p/�//�/�/�/�/�/  ?׿�/6?H?Z?l?~? �?�/�?�?�?�?�?O �?2ODOVOhOzO�O�O -O�O�O�O�O
__�O @_R_d_v_�_�_)_�_ �_�_�_oo*o�_No `oro�o�o�o7o�o�o �o&�oJ\n ����E��� �"�4��X�j�|��� ����A�֏����� 0�B�яf�x������� ��O������,�>��<L������u�����q���ͯ��,������"�	� F�X�?�|�c������� ֿ������0��T� f�Mϊ�qϮϕ����� �����,�>�?b�t� �ߘߪ߼�˟����� �(�:�L���p��� �����Y��� ��$� 6�H���l�~������� ����g��� 2D V��z����� c�
.@Rd �������q //*/</N/`/��/ �/�/�/�/�/�//? &?8?J?\?n?�/�?�? �?�?�?�?{?O"O4O FOXOjO|OSߠO�O�O �O�O�OO_0_B_T_ f_x_�__�_�_�_�_ �_o�_,o>oPoboto �oo�o�o�o�o�o �o:L^p�� #���� ��� 6�H�Z�l�~�����1� Ə؏���� ���D� V�h�z�����-�ԟ ���
��.���R�d� v�������;�Я��� ��*���N�`�r���Ж������@���>�@������ 	��+�=��,)�n� !ߒ�y϶��ϯ����� �"�	�F�-�j�|�c� �߇����߽������ �B�T�;�x�_��� �O��������,�;� P�b�t���������K� ����(:��^ p����G��  $6H�l~ ����U��/  /2/D/�h/z/�/�/ �/�/�/c/�/
??.? @?R?�/v?�?�?�?�? �?_?�?OO*O<ONO `O�?�O�O�O�O�O�O mO__&_8_J_\_�O �_�_�_�_�_�_�_�� o"o4oFoXojoq_�o �o�o�o�o�o�o�o 0BTfx�� ������,�>� P�b�t��������Ώ ������(�:�L�^� p��������ʟܟ�  ����6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z����� -�¿Կ���
�ϫ� @�R�d�vψϚ�)Ͼπ��������*�`�,��`���U�g�y�Qߛ߭߇�,���ߑ����&�8� �\�C���y��� ���������4�F�-� j�Q���u��������� ���_BTfx �������� ,�Pbt�� �9���//(/ �L/^/p/�/�/�/�/ G/�/�/ ??$?6?�/ Z?l?~?�?�?�?C?�? �?�?O O2ODO�?hO zO�O�O�O�OQO�O�O 
__._@_�Od_v_�_ �_�_�_�___�_oo *o<oNo�_ro�o�o�o �o�o[o�o&8 J\3����� ��o��"�4�F�X� j��������ď֏� w���0�B�T�f��� ��������ҟ����� �,�>�P�b�t���� ����ί�򯁯�(� :�L�^�p�������� ʿܿ� Ϗ�$�6�H� Z�l�~�Ϣϴ����� ����ߝ�2�D�V�h� zߌ�߰��������� 
��.�@�R�d�v�ﴚ�qp���qp���������������,	N�r� Y������������� ��&J\C�g �������" 4X?|�m� ����/�0/B/ T/f/x/�/�/+/�/�/ �/�/??�/>?P?b? t?�?�?'?�?�?�?�? OO(O�?LO^OpO�O �O�O5O�O�O�O __ $_�OH_Z_l_~_�_�_ �_C_�_�_�_o o2o �_Vohozo�o�o�o?o �o�o�o
.@�o dv����M� ���*�<��`�r� ��������̏���� �&�8�J�Q�n����� ����ȟڟi����"� 4�F�X��|������� į֯e�����0�B� T�f�����������ҿ �s���,�>�P�b� �ϘϪϼ������� ���(�:�L�^�p��� �ߦ߸�������}�� $�6�H�Z�l�~��� ����������� �2� D�V�h�z�	��������������
�}�����5@GY1{�g,y �q���< #`rY�}�� ���/&//J/1/ n/U/�/�/�/�/�/�/ �/ݏ"?4?F?X?j?|? ���?�?�?�?�?�?O �?0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�_�_'_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o $�oHZl ~��1���� � ��D�V�h�z��� ����?�ԏ���
�� .���R�d�v������� ;�П�����*�<� ?`�r����������� ޯ���&�8�J�ٯ n���������ȿW�� ���"�4�F�տj�|� �Ϡϲ�����e���� �0�B�T���xߊߜ� ������a�����,� >�P�b��߆���� ����o���(�:�L� ^�������������� ��}�$6HZl ��������y  2DVhzQ��|�Q�����������,�/./�/R/9/v/ �/o/�/�/�/�/�/? �/*?<?#?`?G?�?�? }?�?�?�?�?OO�? 8OO\OnOM��O�O�O �O�O�O�_"_4_F_ X_j_|__�_�_�_�_ �_�_�_o0oBoTofo xoo�o�o�o�o�o�o �o,>Pbt� ������� (�:�L�^�p�����#� ��ʏ܏� ����6� H�Z�l�~������Ɵ ؟���� ���D�V� h�z�����-�¯ԯ� ��
����@�R�d�v� �������Oп���� �*�1�N�`�rτϖ� �Ϻ�I�������&� 8���\�n߀ߒߤ߶� E��������"�4�F� ��j�|������S� ������0�B���f� x�����������a��� ,>P��t� ����]� (:L^���� ���k //$/6/ H/Z/�~/�/�/�/�/h�/�/���+������?'?9=?[?m?G6,YO�?QO �?�?�?�?�?OO@O RO9OvO]O�O�O�O�O �O�O_�O*__N_5_ r_�_k_�_�_�_�_�� oo&o8oJo\ok/�o �o�o�o�o�o�o{o "4FXj�o�� ����w��0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� ����(�:�L�^�p� �������ʯܯ� � ��$�6�H�Z�l�~��� ���ƿؿ���ϝ� 2�D�V�h�zό�ϰ� ��������
���_@� R�d�v߈ߚߡϾ��� ������*��N�`� r����7������� ��&���J�\�n��� ������E������� "4��Xj|�� �A���0 B�fx���� O��//,/>/� b/t/�/�/�/�/�/]/ �/??(?:?L?�/p? �?�?�?�?�?Y?�? O�O$O6OHOZO�$U�I_INUSER  ���{A��  �[O_O_MENH�IST 1L{E�  (� �@��(/S�OFTPART/�GENLINK?�current=�menupage?,153,1�O_�_1_C_�'�O�N7�1�@BARRA_ESTEIRA�O��_�_�_�3)X_�Ee�dit�BMAIN>�PLACE0�_o`.o@o�_�_�K27op�o�o�o�o �9`o~�^COLOCA�@�SA_IRVIS�IOa/AS�s� �osm936�����dv�A48,2�%�7�I�[� ���O����Ǐُ�3���0�A����"� 4�F�X�j�m������� ��ȟڟ�{��"�4� F�X�j���������į ֯�w���0�B�T� f�x��������ҿ� �����,�>�P�b�t� ϘϪϼ�������� �(�:�L�^�p߂߅� #߸������� ��� 6�H�Z�l�~���� ������������D� V�h�z�����-����� ����
��@Rd v��);��� *�N`r� ������// &/8/�\/n/�/�/�/ �/E/�/�/�/?"?4? F?�/j?|?�?�?�?�? S?�?�?OO0OBO�? fOxO�O�O�O�O�OaO �O__,_>_P_;t_ �_�_�_�_�_�_�Oo o(o:oLo^o�_�o�o �o�o�o�oko $ 6HZl�o��� ���y� �2�D� V�h��������ԏ ������.�@�R�d��v�aX�$UI_P�ANEDATA �1N������  	��}/frh/g�ui��dev0.�stm ?_wi�dth=0&_h�eight=10�ԐÐice=TP�&_lines=�15&_colu�mns=4Ԑfo�nt=24&_p�age=whol�eÐ��\V)prsim#�L�  }O��s���������ͯ ) ϯ�گ���;�M�4� q�X�������˿������%�\V���    � �]���cgtp/flexÐ(Ǒ̟ޛ2�3t����1
�doubÐ2/��ual����_� �"�4�F�X�j�ώ� u߲��߫������� �B�)�f�M�������3� D�  �������*� <�N�`�����Ϩ��� ������i�&8 \C��y��� ���4Xj���������� �� /S$/��H/Z/ l/~/�/�/	/�/�/�/ �/�/ ?2??V?=?z? a?�?�?�?�?�?�?
O }�@OROdOvO�O�O �?�O1/�O�O__*_ <_N_�Or_Y_�_}_�_ �_�_�_�_o&ooJo 1ono�ogo�oO)O�o �o�o"4�oXj �O������O ��0�B�)�f�M��� �����������ݏ� �>��o�o������� ��Ο��3��w(�:� L�^�p���韦����� ܯï ����6��Z� A�~���w�����ؿ� ]�o� �2�D�V�h�z� Ϳ�����������
� �.ߕ�R�9�v�]ߚ� �ߓ��߷������*��N�`�G����	��������������"�) ��G���6�s������� ����4������� K2oV���� ����#������$UI_POSTYPE  ��� 	 �/�UQUICKMEN  d�s�WREST�ORE 1O��  �	�� /#���m+/T/f/x/�/�/?/ �/�/�/�/?�/,?>? P?b?t?/�?�?�?? �?�?OO(O�?LO^O pO�O�O�OIO�O�O�O  __�?_1_C_�O~_ �_�_�_�_i_�_�_o  o2o�_Vohozo�o�o I_So�o�oAo�o. @Rd���� �s���*�<��o I�[�m������̏ޏ �����&�8�J�\�n���������ȟڟ�S�CRE�?��u1sc��u2�3�4�5*�6�7�8��wTAT`� �<�MUSER������ks���3��4���5��6��7��8���UNDO_CFG Pd����U�PDX�����None���_INFO 1Q�5<��0%��W� ��E���i�������� �տ���:�L�/�p����eϦύ)�OFF?SET Td@���{������	�� -�Z�Q�cߐ߇ߙ��� �������� ��)�V� M�_�q�۹������
���t��)�WO_RK U4������A�S��ψ�UFR?AME  ����&�RTOL_AB�RT��$���ENB�����GRP 1V���Cz  A���+=O@as�����U�������MSK  h�<���N��%4���%��)��_EV�N�����>�2�W��
 h���UEV��!td�:\event_�user\-�C�7���}�F��S�P��spot�weld�!CA6����! �Z/�/:'�H/~/l/ �/�/�/�/-?�/Q?�/ ? ?�?D?�?h?z?�? O�?)O�?�?OqO`O �O@ORO�OvO�O_�O��O7_�O[__Z]Wf+�2X����8V_�_�_ �_�_o�_,o >oobotoOo�o�o�o �o�o�o�o:L�'p�]�����$VARS_CO�NFI�Y�� F�P{���|CCRG�\��>�{�ut�D� BH� Ypk�a�C�� ���}�?���C,&Q=���ͩ�A �MRv2b���	�}�	��@�%1:� SC130EFG2 *����{����Y�X� �5}������A@k�C�F� w�Q�[���|�@���������T��ā�\�ϟ �\� B���;�e�@� ǟ`�����S�����̯ ���ۯ�&�}��\��G�Y���E���ȿ�TCC�c
���������pGF�pgd���-�23456789017�0?��ׁ$���4�v�@Nm�� ��϶�BW������i�}�:�o=LA�څ�6�@�6� ͿZ���i�7����(��W���-�]�X�jĈ� �ߕϳϹ�������� �%�7�I�r�m�ߨ� �ߵ����������8� 3�E�W������}��� ����������/�A��S�e�w��MODE���t �RSL�T e�|k�%" zς��;�1��d���`��SELE�C��c��	IA�_WO�Pf �� W,	�	������G�P� �����RTS�YNCSE� ���$�	#WINURLg ?*ـ�;�\/n/�/�/�/�/�uI�SIONTMOU8���A# ��%��gSۣ�Sۥ�P�� FR:�\�#\DATA\��/ �� M�C6LOG?  � UD16EX�@?\�' B@� ���2T1  �abriel_Fariak?P5�?�?������ n6  ���GV�2\�� -��5�� �  ��Z�@U0>58TRAINj?��4*B{Rd_Cp��D #`{2��'$t�"��h#� (� kI�Mw��O�O�O�O�O 1__U_C_]_g_y_�_��_�_�(STA� i���@��o0oI:$�obo�%_GE�jv#��~@ �
��\��btgHOMIN��kSۮ��`�P2,,��CWǖB�veJMPERR {2l#�
  Qo I:��"�4Fwj |����������&%S_g0REr�m�^۴LEXd�n�1-ehoV�MPHASE  ��e׃BޱOF�F _ENB  ��$VP2�$o/Sۯ��x�c C;�@ �@�;����?s33'D*AA ��]� ��0ޱ�`r}�XC��܅���p\A-۟E �� ����#�5������� ������}�������� ��c�X���A����� ϯ�+��߿��M� B�q���xϊϹ���� ��������7�I�;�m� b�)ߣ�Eߓߡ߳��� ��3���W�L�{ߍ� �ߑ���������� /�$�6�e�W���c�y� ������������� O���?M_q��� ����'9�= 7Is����� �/m/%/3/E/�s�TD_FILTuE�`s�k �x2�`����/�/�/�/ �/	??-???Q?�6�/ ~?�?�?�?�?�?�?�?�O OoiSHIFTMENU 1t}<5�%5�~O)�\O �O�O�O�O�O�O�O'_ �O_6_o_F_X_�_|_��_�_�_	LIV�E/SNAP�S?vsfliv���_��z`ION �ҀU
`bmenu &o+o�_�o�oV"<E�uz��4IMO�v����zq�WAIT�DINEND  a�ec��b�fOKوNOUT�hSD�yTIMdu��o|G�}#�{C�z�b�z�xRELE���ڋxTM�{�d=��c_ACT`و���x_DATA �wz���%  E�GA_BARRA�_ESTEIRAx�o6Ex�RDIS
`~E��$XVR�a�x�n�$ZAB�C_GRP 1yvz��� ,��2̏.MZD��CSKCH�`z���aP@��h@�IP�b{'���şן�[��MPCF_G 1|'���0�r�8�d�� �}'��p�s�� 	(���  �<l0  ���  ���5��>����?��5��`��?5��U��ģ�C�Tp��1V��>w�@3>�?|��/�Q��6 �`��@Q�>���`������˯ݯ� ���o���w����� /�C3�����"��3�� ˿ݸĸ��	��1�@?�i���'�9�0?��Q��	��`~����_�CYLIND~!�� Р ,(  *.�?ݧ+�0h�Oߌ�s� ���� ����(�	�x�-��&� c�߇�������j� P����)��~�_�q���� �2�'��� �&�����������&��I��cA����SPHERE 2������� ���A�T/A�� e����� �/N`=/�a/H/�Z/�/��/�/�/�ZZ� ��f