��   K�A��*SYST�EM*��V9.3�044 1/9�/2020 A� 	  ����CELL_GRP�_T   � �$'FRAME� $MOU�NT_LOCCC�F_METHOD�  $CPY�_SRC_IDX�_PLATFRM�_OFSCtDI�M_ $BASE{ FSETC���AUX_ORDER   ��XYZ_MAP ��� �LE�NGTH�TTC?H_GP_M~ a �AUTORAIL�_0��$$CL�ASS  �S����D��DVERSION  VIRTUAL�-9LOOR 8G��DD<x$�?������k,  �1 <DwX<� y�����C�@����	/��Z �Zm//�/_/�/�/�/$ �/�/	?�';�$MNU>A�\"�  <�:�;"ſ����ZOq?��:�;Uz�m��:n��Z#�o0��ď\�C��/�õ���0�?/ �?'�?�?�?�?�?!O O)OWO=OOO�OsO�O �O�O�O�O_�O_A_�'_�;5NUM  ������92TO{OLC?\ 
Y7 %/U_&2 7_�_	o1_ o?o%o7oYo�omo�o �o�o�o�o�o�o; !CqWy��� ���Z�Vy�Wy