��   �;�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_CPC�_T 4 $�COMMENT �$ENAB�LE  $M�ODJGRP_N�UMKL\  $UFRM\~] _VTX M ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�? �ELAY_T�IMJSPEED�_CTRLKOV�R_LIM? p JD� L��0�UTOO�i��O���&S. � 18J\TC�u
 !���\�� jY0  �� �CHG_S{IZ�$AP!��E�DIS�]$!�C_+{#s%O#)J�p 	]$Jd#�  �&s"�"{#�)�$�'��_SEEXPA�N#N�iGST�AT/ DF�P_BASE �$0K$4!,� .6_V7>H73h}J- � }܏\AXS\UP�LW�7���9a7r �< w? �?�?��?�?�//�	7ELEM/ �T �&B.2NO0�G]@%CNHA�DF#~� $DATA)qhe0  P�J�@ 2 
:&P5 �� 1�U*n   _VS iSZbRj0jR(�VyT�(�R%S{TROBOT�X�SARo�U~�V$CUR_���RjSETU4"	� �bAISP_M�GN�INP_ASSe#�PB!� `C iH�77`e�.fXc1��CONFIG_wCHK`E_PO* �}dSHRST�gM�^#/eOTHERRBT�j_G]�R�d�Tv �ku�c��&T1r
0R HLH�d� 0  lt<Ne'AVRFYhH^t�5�1�� ��W�_As$R��dSPH/ (G%Q�Qt�Q3wBOX/ 8�@F!�F!��G �r{�sjTUI}Ri@  ,��F�pER%@2 {$�p L�k_SF�!�ZN/� 0 IF�(@�p��Z_�0�_p�0wu0  @�Q�7yv	
��
�$$�CL`  �S�����Q��Q��VERSION���  0���IRTUAL����' 2 �Q?  �p�J��&@>�m��`��������������Ғd��Cz  0����A���l��� ������Ɵۯ����  �2�D�F�h�}����� ԯſ�����
��.� @�R�d�fϋϚ����� п���ώ��*�<�N� 	�rχߖϨ�b��Ͼ� ����&�8�^�\�n� ���߶�������� �"�4�F�X�m�|�� ����������� 0�B�h�Vx������ ������,> Pbw����� ��//(:L� `/��/����/� ??$/6/H/Z/l/�? �/�?�/�/�?�/�?O #O2?D?V?h?jO�?�O �?�?�?�O�O__.O @OROdOvO�O�_�_�O �O�_�O	oo�_<_N_ `_r_-o�_�o�_�_�o �_�o)8oJo\o�o �o�o�2�o�o��o �%�4FXj|�� ����������!� 3�B�T�f���z����� ��ҏ�����/�>� P�b�t���������Ο ������+�=�L�^� p��������ʯܯ� ��'�9�H�Z�l�~� ���ϴ���ؿ���� #�5�G�V�h�zόώ� ������������1� C�R�d�v߈ߚ߬߮� ������	��-�?��� `�r���Q������� ����;M\�n� ���������V���� "7IXj|� ������� /E/W/fx���/ ��/��/?,/A? S?b/t/�/�/�/�?�/ �?�/?O(?=OOOaO p?�?�?:O�O�?�O�?  OO'_6OK_]_lO~O �O�O�O�_�O�_�O_ #o2_GoYokoz_�_�_ �_�o�_�o�_
o@o1  Ugvo�o�o�o�o �o��-�<Q� c������u�� ���Ώ8�*�_�q��������ʏȏڋ�$�DCSS_CSC� 2���Q  P����:�܉d
�k�.� ��R���v�ׯ���� Я1���U��y�<��� `���ӿ�������޿ ?��c�u�8ϙ�\Ͻ� ���Ϥ������;��� _�"߃�Fߧ�j߷��� �����%���I��m� 0���f�������~�GRP 2��' ����	ҟS� >�w�b����������� ����=(aL �p������  K6oZ� ~������/ 5/ /Y/D/}/h/�/�/ �/�/�/�/?�/
?C? .?g?R?�?�?�?z?�? �?�?�?O-OOQO<O uO�O�OdO�O�O�O�O _�O_;_&___q_�_ N_�_�_�_�_�_�_�_�%ooIo��_GST�AT 2��%�ߜ< �4���Z�a?�  5O+�ӿ�`�`S�d�Ҵ��aD���:�,DG�	���8`<�e�a܉�e䁠dZCއ���o��c)��}�a�l9E�D�` �cD�`OuW�a\q�`]�`9���DH:�z��c�iD|�/:���`�xN `y���o�o�y��<� N���0�z���f��� Љ�o/g��+k�y �.� �&�H�v�\�~����� ���ȟڟ��*���Z� l���x���|���د� ��.��B��J�0�B� d���x���ȿ������ ����F�H��Ϻ� tϾ��Ϫ������� <���$�r߄�ߨߺ� �ߦ������&�8�� \�n�H�Z������ �����"����X�j� `ߎ���:��������� ��BT.`� dv����� >*t�|�� �V��/�(/:/ /F/p/J/\/�/�/�/ �/�/�/�/$?�/?Z? l?F?�?�?|?�?�?� �?O O�?DOVO0OBO �O�OxO�O�O�O�O
_ �O�O@_R_,_v_�_b_ �_�_�_�_�_o�?*o <o�_HoroLo^o�o�o �o�o�o�o�o&  \nH��~�� ���"�o*�X�� D�����z�ď֏��� ����B�T�.�x��� d������������� ,�>��J�t�.�\��� ��V���̯ޯ(�:� �^�p�J��������� ܿ�ȿ�$���H�Z� 4�FϐϢϘ�����r� �������D�V�0�z� ��fߘ��ߜ߮���
� ��.�@��L�v�P�b� �����������*� <��`�r�L�~����� ��������& 2 \6H��~�� �����FX� |�hz���� /�0/B//./x/�/ d/�/�/�/�/�/�/�/ ,?>?4b?t??�?�? �?�?�?�?�?O(OO 4O^O8OJO�O�O�O�O �O�O�O_�O�OH_Z_ P?b_�_*_|_�_�_�_ �_o�_oDoo0ozo �ofo�o�o�o�o�o�o �o.@dvP� �f_�����*� ��`�r�L������� ̏ޏ��ʏ�&� �J� \�6�����l�~�ȟڟ �������F� �2� |���h���į��Я�� ԯ�0�B��f�x�R� �������������� ,�ƿ�b�t�NϘϪ� �϶��Ϻ����(�� L�^�8�jߔ�n߀��� �߶� �����H�� 0�~��*������ �����2�D��h�z� T�f������������� .dvl� �F����* N`:l�p� ���//� /J/ $/6/�/�/��/�/b/ �/�/?�/4?F? ?R? |?V?h?�?�?�?�?�? �?O0O
OOfOxORO �O�O�O�O�O�/�O_ ,_�OP_b_<_N_�_�_ �_�_�_�_oo�_o Lo^o8o�o�ono�o�o �o�o _6H�o T~Xj���� ���2���h�z� T������������ҏ �.�$6�d���P��� ����П⟼���� �N�`�:�����p��� ̯�������8�J��@��$DCSS_�JPC 2@��Q ( D1����������� ��ۿ�������� Y�(�g�Lϡ�p��ϔ� �ϸ����1� ��g� 6�H�Z߯�~��ߢ��� �����?�� �u�D� V�h��������� )���M��.�p���d� v�����������7 [*N�r� ����!�/ i8�\���� ���//�/"/w/ F/�/j/�/�/�/�/? �/�/=???0?�?T? �?x?�?�?�?�?O�? �?8O]O,O>O�ObOtO �O�O�O�O�O#_�OG_ _k_:_L_�_p_�_�_��_�_�_ch�Sq��u�L�_Uooyo}`d Do�oho�o�o�o�o �o1�oUy@R d������� ?��c�*���N���r� ����󏺏̏ޏ��M� �q�8���\�����ݟ ���ȟ%�����Y� �F���j�ǯ��믲� �֯3���W��e�B� ��f�x���������� �A��e�,ω�Pϭ� t��ϘϪϼ��+��� O��s�:ߗ�^߻߂� �ߦ�������K�� $�6�H��l������ �����5���Y� �}� D�V�h����������� ��C
g.�R �v������ �Qu<�`�����/�&dMO�DEL 23ksx�O(
 <O$}c (  O&z(�/g/y/�/�/�/ �/�/�/�/D??-?z? Q?c?u?�?�?�?�?�? �?.OOO)O;OMO_O �_�OY/�O�O_�O�O <__%_7_�_[_m_�_ �_�_�_�_�_�_8oo !onoEoWo�o{o�o�o �o�o�o�O�O�O�o |�oew���� ��0���+�=�O� a�������䏻�͏ߏ ���b�9�K���3 Es����m�۟��� �#�p�G�Y���}��� ����ůׯ$����Z� 1�C�U�g�y���ؿ�� ��ϩ������h�� Q�cϰχϙ��Ͻ��� �����d�;�Mߚ� q߃��ߧ߹������ �N�%�7���1�C� q��Y�����&���� \�3�E�W�i�{����� ��������/ A�ew���� �������=O �s������ �/P/'/9/�/]/o/ �/�/�/�/?�/�/:? ?#?5?�?/]?o? �?�?�?O�?�?HOO 1OCO�OgOyO�O�O�O �O�O�O�OD__-_z_ Q_c_�_�_�_�_�?
o �?�_�_Ro)o;o�o_o qo�o�o�o�o�o�o <%7I[m� �������� !��_��oI�[�ȏ�� ����Տ�����/� |�S�e����������� џ�0���f�=�O� a�s�����m������� ѯ>��'�t�K�]�o� �������ɿۿ(��� �#�p�G�YϦ�}Ϗ� �ϳ�����$����� ���5�Gߴ�/ߝ߯� ������2�	��h�?� Q�c�u�������� �����)�;�M��� q�����k�}߫���* ��%7I[� ������� \3E�i{�� ��/��F/���� !/3/�//�/�/�/�/ �/?�/?T?+?=?O? �?s?�?�?�?�?O�? �?OPO'O9O�O]OoO �OW/i/{/�O�O�O�O _^_5_G_�_k_}_�_ �_�_�_o�_�_Hoo 1oCoUogoyo�o�o�o �o�o�o�o�OV�O 1u����
� ����)�;���_� q���������ˏݏ� <��%�r�I�[�m�����$DCSS_P�STAT ����ӑQ?    �� � (�+��4O���t� r�Ԑ@���������é���ӕ௎�կ�ĔSE�TUP 	әBȖ�ãá8�R��ͬs�b���������T?1SC 2
+���ƱCzƳ���;صCP R�D�DLj�|�>�� ���ϓ��������0� B�T�#�xߊ�Yߛ��� �ߡ�������>�P� b�1����y����� ����(���L�^�p� ?��������������� ��$6Zl~� Vϫ�D��� );Mq��d ����//�7/ I/[/*//�/�/r/�/ �/�/�/?!?�/?W? i?8?�?�?�?�?�?�? �?�?O/OAOOeOwO FO�O�O�O��O�O_ �O+_=_O__s_�_�_ f_�_�_�_�_oo�_ 9oKo]o,o�o�o�oto �o�o�o�o#�oG Yk:����� ����1� ��g� y�H������������ 	��O-�?�Q�؏u��� ��h���ϟ����� �;�M�_�.������� v�˯ݯ�����%��� I�[�m�<��������� ٿ���̿!�3��W� i�{�Jϟϱ��ϒ��� �����/�A�S�"�w� ���j߿��ߠ���� ���=�O�a�0��� ��x��������'� ��K�]�o�>������� ����������#5 Yk}L���� ���1Cg y�Z߯��Z� 	//�?/Q/c/2/�/ �/h/z/�/�/�/?? )?�/M?_?q?@?�?�? �?�?�?�?�?O%O7O O[OmOONO�O�O�O �O�O�O�O�O3_E__ i_{_�_\_�_�_�_� �_oo�_AoSoeo4o �o�ojo�o�o�o�o +�oOasB� �x�����'� 9��]�o���P����� ɏ�����Ώ#�5�G� �k�}���^���şן �������_C�U�ܟ 6�����l���ӯ寴� 	��-���Q�c�u�D� ����z�Ͽ��¿� )�;�
�_�qσ�Rϧ� �ψϚ������%�7� I��m�ߑ�`ߵ��� �ߨ������3�E�W��c��$DCSS_�TCPMAP  ������Q @ c��c�c�c����c�c�c�c�	�c�
c�c�c��c�c�/�  �c�c�c�c�*c�c�c�.�c�Uc�c�c�c�Uc�c� c�!c�U"c�#c�$c�%c�U&c�'c�(c�)c�U*c�+c�,c�-c�U.c�/c�0c�1c�U2c�3c�4c�5c�U6c�7c�8c�9c�U:c�;c�<c�=c��>c�?c�@u�UI�RO 2��������������� ,>Pbt� ������	��-��Qcu� ������// )/;/M/_/q/�/�/ 2�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O�/3O�/WO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_��_�_&O�_q�UIZ�N 2��	 ����� oo$o*��_ Rodovo9o�o�o�o�o �o�o�o*<N r��Y���� ��&�8��\�n�=� ������ȏ������ ߏ4�F�X��|����� o�ğ֟蟫���0� ��T�f�x�;�M�������������_x�UF�RM R�����81�^�p�/�� ��ʿܿ�� ���6� H�#�l�~�YϢϴϏ� �������� �2�I�V� h�ߌߞ�y����߯� ��
���.�@��d�v� Q����������� �*�A�N�`������ q����������� 8J%n�[�� ����"9�F X�|�i��� ��/�0/B//f/ x/S/�/�/�/�/�/�/ ??1(?P?b?=?�? �?s?�?�?�?�?O�? (O:OO^OpOKO�O�O �O�O�O�O __)?;? H_Z_�O~_�_k_�_�_ �_�_�_�_ o2ooVo hoCo�o�oyo�o�o�o �o
3_@R�ov �c������ �*��;�`�r�M��� ����̏ޏ����+ 8�J��n���[����� ��ǟ���ٟ"�4�� X�j�E�����{�į֯ ������