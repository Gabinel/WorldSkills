��  	^��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ��!PCOUPLE�,   $�!PPV1CES C G�1�!�� A> �1	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q�RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Nb_OPT�2 �� ELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1� UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t���MO� �sE 	� [M�s��2�wREV�BILF��1XI� %�R 7 � OD}`j��$NO`M��!b�x�/��"u�� ����4AX��@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC���a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���OR BIGALwLOW� (KtD2�2�@VAR5�0d!�AB e`BL[@S � ,KJqM�H`9S�pZ@M_O]z�ޗ�CFd �X�0GR@��M�NFLI���;@UIRE�84�"� �SWIT=$/0_N�o`S�"CF_�G�� �0WAR�NMxp�d�%`LI��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqS��� X�r$ORIأ.&ӧRT�`_S�Fg�0CHGV0I��p�T��PA�I"��T�2@��K�� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8��9�4��x@�2� @� TRQ��$�%f��ր����_U袰����Oc <� ����Ȩ3�2���LLECM�-�MULTIV4�"$��Av
2FS�ILDD��
1g�Oz@T_1b � 4� STY 2�b4�=@�)24�p�e`DԼ� |9 $��.p��6�I`�L* \�TO��E��EXT���ї��B�ю�22�0D��@��1b.'�б9�G�Q� �"Q� /%�a��X�%�?s��EӂU� Sҟ�;A�Ɨ�M8�� � CՋO�! L�0a�� �X׻pAβ$JOB`B����f���IGO�" dӀ�����X�@-'x���G�ҧ3AC�`\��b# tӀF� f�CNG�AiBA�  ϑ��!���/1��À�0����R0P/p����$
�|��BqhF]�
2J]�_RN���C`J`�e�J
?�D/5C�	�ӧ���@{ ��Rd%� �����ȯ�qGӨg@�NHANC��$LG5��a2qӐ��ـ�B�A�p��z�aR���1��Ex�>$FDB��ERA�cEAZt@�ELT���в`WFCT���F�L�`��SM� �I� lA�f��f��&��5�5����S[�g���M�0��`���#HK��AEs@͐���W��N���1CpXY#ZW�`�����&�	�ѯ���&�2�!S�WAq�"��'p�ST�D_C�t�!W��U+STڒU�()�0U�0�%E�1�!�_�Up�q�) \�1UM)1ORzs>2p;�d��`O< RSY�G� �qd5Up��H`G���{@0A%0PXW�ORK�*Ѱ$�SKP_�pQ��0D�B�TR�p + �C �`����`m�fU DJ�dp�_C"�0;b�3 �7PL:c�a��tő��D�AGQ 92���Q�PV.�P�O�B��,�2&1P	R'��
$0Ja9��g- /�q$r�w$Zz��L{II.�O�����/�O^z�PC�0�O��DENEM�c� 11�O�C\@RE4��B2H $C)bo-$L>S.${C8ނ�O[INE�]13_D!V`ROyp� ������q�S=�z0�V�PA���Rp`RN\�R�MMR(�U��vI�CRmPEWM0^�SIGNZ�A����U�a/$P�-�0$P�s�	1`�`-ds�1`DIp �-�hTTQ/b�GO_AW���h0ؑH!�0CSd��.�CYO�3���P1�}��avIG2�j2vN�}��K�c�c~O�4 P $���RB���PI�gP�KwqBY��p(wT�=A�dHNDG�AG5 H4��!wE��~%�$DSBLI󠌳us�fm0���cL�۱6Url0]��xFB�|�FExQ>��rP�d�c5��7D�i�8Z!���MCS��pPl4&��ra"H�W� K�����L����0�aoSLAVQ8��INP^�(v]����a���9P + �S � � ~�0 �0��FI2����烤�-1�-1Wr��NT�V��Vݑ��SKI�TE`5g�@�$�Z!J�#@#_�@j��SAFT�a|�_S}V��EXCLU��*T0pD\0Lr��Y�t��Y�HI_V< b"PPLY@6�pёS���ӓ_MLs��T0$VRFY_t�3ђM��IOCц[�C_��2��O�p֕LS� |rLD4�$AW��c�о0P��5,��`)�AU��NFzv���e���`s�:1CHD��up�����ЛAFI�CPr�T�$A�r5�_�q :�P�0T��� z� ��d_N��c� I;���T��� ���E�O��SGN��<A 
$ �P�QdQ�� o�9���#��2s��2��ANNUN�@�����e IT0`5�˹`ȱ�к�"2EFi0uI�B=v�$F��4 OT�P��LDj��NB2Ab�IA�M�pN�I�B>��Z��\�Aܼ�x�DAYC3LOCADtADS�MC5IA��EFF_AX�I�r?P7AU#O����C�0_RTRQ���@ DWp/P��Q
�"��E|`�ø����?���� �������AMPE�� A\�6���6�Jc���DU�P����2CAeB��B�PNSH�6��ID��WR �3�4\�VwV_2�������DI���$Cߜ 1$V�PSEs�TWp��M��ژ$@dE_��J�VmE�� SW�@��a ��������@ f��OH��O�PP�&K�IR1B�0�� Lӥ��R�!氃�}#}�@��}�vs��B��x���`��RQDWl�3MS} ��AXR��J�LIFE�0��SA�N�(�ȱ��C�wǳCH �raN*�z�R��ȱO�V 4�HEw�SOUPPO�0{q�"�0_��y�W�_���ma��Z��W��H!��0�ȱfrq"XZerAV��Y2C_PT�0D�P��N���ȱJ�� d�_��!H���C�T�$D `�`C�ACHR����SI�ZN�z�b� SU7FFI�����0�N�AD��MC6IA"2M�v vE 8԰KE�YIMAG�STM RQ\�Q����2W��OCVIE)�01F��"�L!�n�ރ?�K 	��D�vG��m@�STM�!i $@q2@q��q��qEMAILq��P��{I�עFAUL�B�H�"�S�3AXy`U�� �P�@DT-P�!I�< $��S�2Г�IT}sBUF@�ށ��d00��	B$tC݄ԡ�3�SAVS%"��: �3�n'��̶PZ$�0P*�tp_ 9%r��)#OT�R��ңP�:@�*��'AXC3	���X z��#_G�
?��DYN_t�J <WpDuA@�uUs�M^�n�Tr��F�P$�P��DIB��E�0-P.��1K�ǐG)!$�&m�jQ`1�m�p�Fyp L (PSVw`�dADM�6�*d�2�Q3Q�M�:P�1��#C	_�P�PK�T @���4�w�R��5��1DS�P�2PCAKIM@`#8C^Aߥ�1��UG0��U ��IP"��3]�Y 7DTH9 �s+B2��T�Q8CHSk3CGBSC/�H PV����J�@�#�DD`��NV���GS�D9 5F F�� 0dC[0�!�QSqC��u�3MER̔>yAFBCMP̓�0�ETa� N�FU��DU�v��PڒCD.I�@� ��PQR-���c�O���`��Rr��T��P,��RC"H��U0�2U�S|� �PH *�QL����a�!cV�b� M�Yd��WfH�Wf��WfP��Wf�Wf7Ti8Ti�9Tj�Vh`j1mj1�zj1�j1�j1�j1��j1�j1�j2�j2T`kmj2zj2�j2�jU2�j2�j2�j2�j�3�j3`j3mkzj3��j3�j3�j3�j3ʻj3�j4�b�EX	T��c�Q22�70K��70QeB0���Un F{DR��RT��V}��"����B�R�EM�Fla��OV�MC�A�TRO�V�DT^ /�MX�>�IN�`�.���INDM�g
y�l0 050G1��8�_(��9D��8�RIV��L����GEARAIO�K��J�N[0호���*���K�Z_MsCM ��F��;UR�RS ,�Q+!�? _�s@?\K��?K�EV��S�mE!oPՂT j��P�!��RI��p�#ETUP2_� U ��#TD�@V�$T��c������1l���C,2V T(j����4)�:%�cV0�PIFI`�V0oP�@`��PT+��QF�LUI\W ���>�UR��>!f�@�"s1�@ ���I�u$��S;�?x���J�0CO� �#VR�T��%�x$SHO8�װ�ASS�@�!8N��@��BG_�s鱀
��zc鱇c鱔cF�ORC�ID�DAkTA��X�FU6�	1`29�2�5E�9 ��wY |��NAV� ���������S��L�$VISIl���SC�$SEq��Ӱ]�V��O��$��PB"�`�gй�$�PO��Ik���FMR2҅Z ߂�P�����0�� �����&��������_�a���IT_�5��T �M��ɟ۝D�GCLFa�DGDMY��LDc���50�H��(�0�M�`^[%�R� T�FS� ]\ P��.�3> 0$EX_.�E�B.�1� 4Pk�/�3g��5g��GQ��] Y����RSW<%O��DEBUG����GR UVSBK�UaPO1)p "�PO6������P��:��MҰLOO�#�SMb�Eb"ۡk�L�_E ^ ~|��TERM7�9_@�&aORIy1<�}`@�I�SM_�0���<�a@�n -��b�@���UP3c�3 -j���^��N����_��G����EL�TO�d2PFIG�e16��ᆠe����`$UFR���$�P��) �Um�OT�6PTA�@��HN;STz0PAT�A� �^PTHJ�Q�PEt_�3��ART{ �����{!�d1REL<�
�1SHFT�Be1d�_��R�P�S}�% ��$��� b���8��sC2SHI� ���UPb u!AYLO �@1&1H�t�ɲdY��U�@ERV_`/}� ���Dz0��q'���
�'�RCs��UAScYMY1�Ue1WJ���E����}��QU�z0&1���~�aPqCL!QORz0�M�� ��&���d�4����c # 1+�H9O#��e �J+�,���POC�����$OP��AAEcFճ�����0��2� R5S�1OU�Cdem�Rb�%�(����e$PWR��IM�%`R_�#���~�we1UD���0|!�y4f��$H�5!^q0ADDR��H)�Gf�11x1 �PR\��2ag H��S\P ���s�5
��5zc�5�ccSEVѧ��PHS�P���h $~�� _�D����ɲ�2PRM�_i�a�HTTPu_�PH2ai (�P�OBJ��x2��$���LEU�04A3`j� � ��yQAB%_z�T�BSp �C�W�KRL'9HITCOU�D갟 ��� ��B����ų� )�� S�S~�RdJQUER�Y_FLA��yQB_WEBSOC��G�HW�a��2ak�0} INCPU{���OEV�A_d\R�4]Q��4]Q�b �IOL]N�l 8��R�ބ�$SL��$�INPUT_��$� �XP�� G�PSLA�� m�P�_�U�T��U��x!IO@F_AS:�n�$L�ZG����92`��S��S1HY��ca<c�k�`UOP�o `(`�a��]�Sd]�Zf�a� P=3� �g�aZf��b�f�1IP_MEܻ�M�p X(`IPx0{�r_NET{�P���"��"vQ��DSP��,@�ްB�G{�B���M�M�q3 l_�TAGa@A#�TI�e
%= 6�l�u� PS�vBU6�IDZмB#�u� �u0a�[r�rV r�Rmz�t�t�PN �6����IRCA�� �s �xI�PCY�0EAKcB���G�]�=3_���R~ ��s�!DAY_�p�xNTVA\��p���R���s��SCAA��CLڑ�qɱ��r��M��t�����N_�� C-� ��r��N�u �R+��#S��aUB�p�q�@��+� 2t !�P\q��M�v��UB�pLABV��6�.��UNI/���h��ITY�c\q�5bR� ��w�Rd�R_U{RLk��$ALЃEN������~�STT_U�� �J4DPM�x�`$;��D��DPR�e\�t�A��d�Qf�J��r�FLP�䂰�
����
�U�JR��y �x@F�X���"��D���$J7@O�$J8ܩ7��������7��ؠ8�ۡAP�HI��Q�+�D�B�J7J8ɲD�L�_KEِ  ��KPLM
� 7z <�XR`RP�ȳWATCH_V�A��L�QFFIE�Lpu3yb�`���{� i�LVU7���C�T
�̶u �LG~��|� !4�?LG_SIZ�D��`���`�FD�I�"���
�9�� 	��#Ä����`�� 9���9��ƪ������_CM:��W���D�AF�����	��$(���"��"�`"�9�.�I!�8��0"�9�"�	�RS��s �  (���L)NС��}�`�@�� W��RO����C��p �L�Ӯ�DAU��E�A#@P�$����GH��"��+`BOO�1�~� CBb70IaTS� >fREbp�5�SCR
ЪCCaD�I=cS# �0RGI,�$Di��V6c�$��$�D+aSfC*bWq�+a���6cJGM��MN3CHS+aFNV���1K��$���UF��n��FWD��HL5�STP��V��Ԑ��,%���RSm�H& �3fCK��6cT ����UA���:ӳ�ְdKc�G�� PO	�P�`�K�����Nq �E]X2gTUI��Ii� 9�>�i��~����ّ� ��:�	؀R�� vQ�NO�ANA+b�!��AI�D��DCS���3�3O
OSy�4!9S-��IGN"����4����b�DEV6��LL�T��s��`���qT$�$@��MR8�zaK�Ag1���	��PXSq�� OS1�2�3��\�9�`� �xK���U4�T�u�AU$ 3���h&ST��`R��Yp� �  _�$E�&C�+�Р@�&�&��9�a� L?PQo��fh'v�#�@97EN#@;4����~Q�_ � @��)@ՃR�J3��M�C��� �x@C�LDP�`N�TRQ�LIґP�~9l4FL Sq�2A�3�D���7�0PLD�5�4�5OR�GV���2��RESERV`T�4lS�4wR�]3��� � a	�5��{4�5SV�Ф~0��	�1YDaFRCLMCoD�?O�Ix�PaA��MDBGa����m�$DEBUGMASTc��~�J��U��T� �uE���q\0FRQ��߇ � ��HR/S_RU�Q1U�yAc���FREQ��'�$� �OVEAR�p4�p6&��P�7EFI�p%�!V�p�A5�R,D� \F��?Q��$U< S�3?6@��PS�q�	JSC��pC|r�S�C�U��A?( 	�zaMISC��� Yd��<!RQo�	@p3TB|��p 3f��@hAXs2[�Cg\lE�XCES�!bM�`����'bs4/1�bSC=  � 	HP�7d_��1hf��k(Zolh\0K����Rݢ�|��EB_ްFLI�C�$B?�QUIR-E��MO&|O6{�V�$AL0M��� @D0-�sp�soB�A#ND�џ�����Ҡ�����sD�ü�INAsUTb��RSMѠ��xYN�"����q$�L�sPSTL���� 4�LOC?&R�IԐ?%EX4�ANqG��Q	QODAU��#`����L�MF�@�qVe)2��58�����FSUP(68��FXi�IGG1� � �6@3���C 3��4�R�"牌  ��� ��`&~���QCTI��鱉`��MY�n�B� t�MDd��Ȓ)r�
}��Az�H8H��}�DIA�~��l�W��}���}�D��)��MO��W@���� �`CU"�VP��Q@�QaO��_�@��� ���G#q��@&�R�D�.�P.�x�4�5�P-�KE�򌰎�-$BYP!�� N�D2�B��~�2_T=X4XTRA
����B�spLO�з����b��/b���Җp���أ�rRR2e��� -С��A�^A d$CALII9`��G��2��RIN� �<$R�*�SW0�DZ��CA;BCx�D_J��-q\�Pq�_J3��
�G1SPް& �PP�B��3����� �Pյ�J�C� BVAO�IyM�@�RCSKP�:������J���RQ��E�+�E�;�=�_A1Z]B�w�EL���AOCMPK� a�Qƴ�RT�A��ҥ1����=`1��ȩ ��Z��SMG��U��D;JG<0SCL|`8�SPH_9�Pe������P'�RTER$Y� �� �_� W1�d A���#�RU�D�I���23U�D�F�v�LW|�VEL~1IN2� ��_BL
�R����Q�J�Ԭ��׽�L�IN8�?Q�`����Ջ������ _` �@���]���b��mֈ`DH|`���a��$V)��sө�$��UQ8�o�$ʖ��`R蓶`�H �$BEL��|W5�_ACCE��� ��A��IRCi_V�p��0NT�Q�i#$PS|`q2L�<���3����m��� ��u���6���6�3��a_���g�m�PU�P��_MG/SD1D��V�8�FWa0V�`��������DE���PPABN�RO�EE}����~0;����A�`���$U�SE_(��PYPC�TR�Y���\A �!YN`A� T����TM�A ����O8��(�INCڔE�����@b��AaENCF�L<��R����>d��INq"I��W���NT�Ӿ�NT2c3_z�8�LO��8�.gPI�p��9��@0c�@8�0��bC��MOSI���b��m�OS�RPERCH#  UeQ;� �K� ��;�D��Ǖ�>HD�l��Aa��L4 ��g� ��;6&QgTRK9�1AYԣ ��af!a�u%j#F���8�a�PMOM�@b@�b�0��/d����#�8��DU
�b�S�_BCKLSH_Ca��%�@vfP\�S�3�!:k=�CLA�LM��A� <�S5C�HK�H���GLRTY"�o��I��1U�9_��k_UM�C�6�C�C��Ѿ33PLMT��_L�0���4���7E�=�0�;�0���5��跰�C ">D�PC���HTp���5C�MC�����CN_b7�N���F�SF���V>G��5�rAa���EvHCAT�>SH ��7�����1�!�ѥ0�ѩ����PA�4�_P�5�#_��m&`��}#�T�5JGx���`�S��OG�GA�TORQU0 ��i�)���r�B����R_W �%f$����d|�e��eIkI(kI��F�^�a�gh����VC"��0�a�e�b1�n��8�o^��fJRK�l�b,�f�DB
�M&�M�p_DL|�"GRVdt|�t���a�H_ף�c9�@zCO1SM{��MxLN�`p{ �ewt|�ry��ryDa�z��|ba�eZkp��aM�Yyq�xYrw�a{�T�HET0��NK2a3��7�v�zpCB<�kCBv�C,�AS=��a�Ddo�|�o�<�SB8|㍂G�GTS�C��iQ��XS��Ê�s$DU}0'��(������Q�_RC*Q+NE�%�K�4��[�Z�+�A/�X�a�?uJxJqLPHMu6�6�S�e���u���u6���vӓ���vX�Vz�V�o�l���V��V��V���VʛV؛V�V��Hz�������Q�����H��HʛH؛H��H��Ok�Oz�OT%���O��O��O��UOʛO؛O�O�v�F6�\����u��m�S�PBALANCE�_�q�LE��H_/�SP�эvv�>�vPFULC�;°#�;«u��1���U�TO_x0�5T1T2|ɼ�2N_1�� �����!=����!�T' Oo���`IN�SEG��ZREV8��Z�DIFP%"�1��m�1�C O!B��C1s�'2�P�j1�dLCHWAR���CAB_Q�%$MECHe��psy��6AXs!P!D��Q�]�q�� 
���Q��n�ROB�CRa�X�ՇBa��C��_{R�T � x ?$WEIGHp )P#$k��PIp6sIF(��LAGa�@BSa��aBIL�G�OD� ]%�ST��%�P��C0&��� P���О�
� ��b�{Q  2�h*�D�EBU6�L.�v���MMY9����N8IS��)P$D.��$���P� � �DO_��A�џ <�����1$bN�B`�X�N�3��_?b  }�OP0 ��� %�0T�� ��1T������TgICK7�K�T1 �%��� ��N�k�'��R0b[ң�[ү���PROMPpE~M� $IR�P�`�0��
 )MAI��`�r_A��
�|!t RpCO�D��FUh 3�ID�_�E�����G_�SUFFD` h;�W
��DO��0����Z��GRA�[� ���[Қ[Ҧ�Q�������H1�_�FI��9�OR�D`� ���36�%B�` �$ZD�TL��~�
��4{ *	�L_NA<����S��DEF_I cS��o��g��q�`��������IS�@�@�.������mD�A��4�A8Bq�Do�(�"$��D�PO��LOCKEIQ}��`������} UM� S������� �#�~���o��& ��f�|Q�S�� ��')5V�P/��f��4���Wd(c5Z#�� �TEN1��� ;�LOM�B_}2�70%�VI]S[pITY%�A�Q}Oa�A_FRIlÌ�30�SI��1 �R����7���73��%�WB�8W�;p�6�`_4I�EAS-��Q�4P.P* 	�64�95�9�6.�ORMULA�_IIQ�GC�� h ��7��C?OEFF_Ou���H�Du�G!Q-�S6����CA=�����}�G�R� � � �$Z ��(�Xe�TMM'ETZ%{�b#_\1�ER��TC$B�࡛  e�LL�" S�M�_SV$�X$Ć6���p�D�� �7RSETU�MEA��b �`&�}��>�Х � �P�� ��@a��a2!D)fX��2!N!/$�RA�Yc��+ ��* ek�2� R�EC#a�MS�K_�+S� P~�1_USER���4ҷdJ��t�`��VE�L\b�`J��b�e[�I�,���MTV�CF}G�a�  ��z�O��NORE���;�r�K�r� �4 c|�3��X�YZ�������� �3p_ERR�ѩ ��PT�5 Szp����`�`��BUFI�NDXOa�uqM�OR+T� H�CUzq;���q+�c<���$���vA�Nb�A���G-R�� � $SI`�@@5 ���`VO(�<#���OBJE.�)��ADJU��+�:�A�YWP��2�Dh�OU�� Su�pa�=��qT�����`��
�DIR����
������GDYN&B�B߅Tp��S�R�1f�`�R��O�PWOR9� ��,��SYSBUH�PaSOP!��r�Q,�U+�
�PZ �bR��PA�`#aT�}�PaOP� UR�F�/ђ��ჀIMAG�q����q�IM�q��I�N4@z���RGOVCRDԁC��`��P���������0#����L�X Bwp��aPMC�_E4�q��NH�M�$�����1��`ԑS�L.��`� ��O�VSL��SX2DEX!�i�2�����A_Ԑ��� Ր��� ����������C��U��xϡ��Ր_ZERqqH��S�a� @@p4좜�OM RI+���
� �2�%�q�*E�L�a��rT~�u��ATUS`��C_T���rm�BIPw�`��"d#��L�4�`� D�l�j�ܰ��k�0����a��XEq�*eŲٲ����	��p�cUPXd��PX��ȗ�����36������PGu��$S�UB_����!_�3�J?MPWAIT���w�LOWMs|�)�E��CVF����z�RX��p��CCҠRց�����IGNR_P�L3�DBTBu�P����BW1 ��&pULH��IGj���I��OTNLN���R��S"�0N��c�PEE�D�r�HADOWu���&p3�Eq�kԀ��I�nSPD�a� L�A��o��M���CUN#�:˗��RఆڣLY)��i�=P�H_PK5u�rRETRIE3�*r���z�����FI8r�� �X���� 2}�pDBGLV��?LOGSIZ,�!KKT��U�SP�DV�n�_TX�EM�@!C�aۡv�_�Rp�L2>IvCHECK
�Oa��P�`�Ѷ�p�鿂LE"�RPPA�A T��a�ms�IP4Ҏѷ�BARC�8Ӱ��E�O� Nr�@ATT�ҖaC�v�0)b!.��UX��梱PLJ t� $�qM1SWITCH�r�QW6�AS3����q�LLB�ѹ�� $BA�`D(#PaBAM�ă��3���J5jp q���6����_KNOWh��ԀU[cAD���P��D�`%	PAYGLOA#a� C_�q�L$�LZIL�!A�a�LCL_�p !�P����a�*��F�	C�P�
("b��@I�R�P�$�r�BU@�qJڢ
�_J��a�qAND�rsb(��F�@A�PL��AL_ ��~���p����0C�\bDHE[b�J3�=Q� T�@PDcCK��PaCO�P�_ALPHa�BaE�q�Aas �
R|�� � �LЮBD_1I
2sD�PAṞ$(%5& #^�TIA4O)5O)6\bMOM�p[#{#�h#{#u#pB��AD�[#�&h#�&u#PUB�R�$�%h#�%u"���r�d�� L$PI֤2� #�aN9�ɡh	9I*;I8;I F3, mq�w6-�w68������s���O�HIG��Oӏň��6�� �������6�3�8���9<����SAMP԰�v�2D�73C����. o�aA�pq��rpD-� zF�� �I  �r����X xEM��H �zCIN�LMC�H�K�D����J
X�D
[*[GAM�M�ESs�_t$G#ET�2�pQ�D��b;
$TIBR�0�]Ijw$HIX`_đH�p�r�VE�p�XA�^�P�VLW�]�V�\�Y@f�V��6&�SC��GCHK���`�I_@���tL�L��Etg�#�t�&siQ ��$� 1�� �I1�RCH_5D����RN��V��bLE���2� x���`�3�MSWFL���MQSCR"�75��L�pD3W�Tv�G �p[ �Ihy��wt�r�;SV�ѾPـ���;w�qGROU��S�_SA�����u�NO�C����p}T �TfL8:�*�r0Xz5g� #DO��AzR ��qEjz�E�8&��6��`�8ˇǅ��� F��L�`�$� � FycYL3��G�@@L��W����%�	���d)����;p��ñM_W�pk�q�� i��b��M����� ��P���:�q�9�-�� M�q 2� �!����$Wݐ`�ANGLF�vݐ�ے�ے �ےu���PN��S(��q�MX��O�L�Za�� ���$� �,aOM�c��!� 3�E�W�R ��b����uL�_x�� |� ���p{)'�h#'�u#�p�T*T�?�n*��wU (�@��r��w ��P��PMON_�QU7@ � 8���QCOU�aY�Q�TH�HO�ҰH�YS4�ES��ҰU�E���r�Ov�� � ��P���U�qRU�N_TOI���O�2�p� P? ŭŞ�qINDEp�� G�RA��h�*�2q�N�E_NOf��ITx�`h���INFO�q����Nˏ�(��ؑO�I��� (�`SLEQ�6���5��Rƹ��OSM`��� 4���ENAB	��PTION(�k�2�����GCF�� �@��J��L#���PRK����,����EDIT�q� ��!�b�K��3�QE�PNU�מ�AUT<�q��COPY�ѭ0(�܍1�pM�QN����^EfPRUT� ���N=�OU��$G� �+��RGADJZ����X_r�I�cP`�W�n�W�WU�PU�pW��3G��RN8_�CYC	���RG�NS����@LG�ORc�NYQ_FREQ�"W�@�6��B��L~ *���U�v#�@�5CRE�PݳS`�IF81Z�NA;A�%&�_G�cSTA�TU��c�MAI�L9BIqʹLA�STq���ELE�M��� �5�FEASI�˂fB^p Qp��1�q��ҭ@�PIs��d��1ձ��s&AB�sE_��0�V��
*	�R�!U��0�0�pSRMS_TR L�`�nY��0�R��R ����#��	�� 2� �CF��D ������@M�8�7�dDOUH��d�N/Ӽ�PR����О��GRIDm��B7ARS�7TY�ؑr�@O� ��� �E_B�!��i)O_�>��� � q����PORHÒ6�S�RVF�)��DI�pT ���0��0��4�Kp�6�7��8���FZR���~
�$VALU9��u������F����� ! ���\�|H�x�AN�sp"X��R������TOTA�L8C<��#PW��I|1�$REGEN�*�"�X_0��噱�&Ƹ�TRE�2�!_S�pE7� �VU�p�f2.�Ex�5ױ���ܸЪ#V_HRDA8��e0�0S_Y�qY����SFpAR��2�� #�IG_SE���O0���_��4C=_]$CMP��BKDE ��0BIUa�ZC�3�QCG!EN�HANC��� �p��X�S�1I#NT��!��F�}��MASKT�P OVRݳP��5ԠG�aF�E#4���B��|;]�PSLG�0
���C��r��Qr���� � SX���!A1UPq�STEQ�P G��� �QEeJ�F<�r	�IL_M��Pso0��TQ���Cr��Y wL�V�[C�]P�_�P�p�SM�YV1V�ZV1�[2	k2�[U3	k3�[4	k4�Z �qk0kr�q.ІfZ�lr;IN�iVIBȐ�T��`���d2�h2�h3*�h3�h4�h4�h����RِS�r���T $MC_F۰�p��L�q�qaE�� M�pIaC>r
 ����!Bo�KEEP_HNADD7q�!yt# �yC��F� �ti8r+P�sO��xt��6qn0�sfG�sREM�r�t�!��u�q��xUB�e�tHPW�D  ysSB�M�A�COLLAAB���  P�!,���cIT��P���NO���FCAL �u}�ڛ ,��FL�IO$SYN0p��M���C�2�� UP_D�LY���
�DEL�Aɀ�!U�Y��AD����AQSKIPNߕ� Ģ�O+�cNT�aM��P_� F��N�E�� )�k17� .�7��6� 6� 6�@& 6�3 6�@ 6�9�O�J2R�������XD T��ؑ����ؑ�D�urؑm�uq��RD�C�!�� ���R"L�R���P�aR�"�8ղ!��RGEY���)�FLG����9�9W��SPC�ç��UM_ؐwS2TH�2N��ː o1� 	�EDi>�� � D;�[H<q�' 2_PC����SIQn���L10_�C��м��A �O�$젘���*� ��R�Q+�)���hѪa��)�b�]��"�2�'�A��t@Ǡ�9�Dr�G��VL1멱1�����10�p_�DS�Q�Q~�5��11��� ljp�q<R�p�]�AT�p,� ��'�R�V�����¼PҞbHOMEH� �2������"Ϡ4�F�X���3���{ύϟϱ�������4�����
��.�@�R�W �5���u�@�ߙ߽߫�����6��������(�:�L� +��7���o��0������ �d�8��������"�4��F���S=�v��  ��0m���p=E�� T͠��L�&��IOtQ	I��:�2Oy�_OP*Bx�"l�j�POWE�a�� ������¾$ 푅y$wDSB!PGNA��Ľ#ĀC��r!��S2;32� ��n���pHPICEUS��#SPE��i!PA�RIT�1�!OPB�e�h"FLOW�0T�R���"�qU�3CU8� J�j!UXT�Ai!>t@ERFAC��p�U� ��SCHN�� tjp3p_� �@w�$�0�0OM��02SAR�7�/@9qUcPDPp
�{�PT���EEX���nPE�FASp B�1M#�# сh@�" �SZ"� �a���qK!  2� �S�~w��	� �$��Bم��c%?#� _�0�J&DSPV&JOG@t0���n�N͐�ۅ���6K�_McIRr!�$�@MT�S�#AP�S�@��� D��S�0� .���@�%�BRKHi���A;XI��  2�C�2A"�A�2?#� BSSOCJ&�pNF5D�0�Y16s�$SV&�pDEG�F�G�PeD�D�B�#OR�7��N^@�6F0�7o OVr%SF�:�0�3�BF�6/�#UFR�A�:TOLCHXǂۅ�POV�En!WE�K�o#�q�2S0령_�0]� @|�T�INVE[ ��OFeSp@C��SWD�1�3D�1R1z��%l0TR���u�E_FD<��!MB_Ck��BB�B�P>����B�AS�y0V�q�R�:�ك2�2G�G�(AM�#�@0jUZB5__M�@/s�g@T$	�)P�>��T$HBK��&�QIO���U:�QPPA�Z�Q�Y�T�U�@U:gBDVC_DB3����P���PK�@/	e�`hZS	e3f@`@Y���?� �1U��d CAB��򒣠�@L��@X��O(PU�X�&SUBCPU�| S1�C��T��C��i�CTv�$HW_C���C��P��fS����p��$�Ud�#4ppAT�TRI|�*r| CY�CԢ{aCAVb�#F�LTR_2_FI���	\c��P�+C{HK+�_SCT�#F_wF_ |�r2z�FS��BrCHA�1��w�q�B$�rRS�D���31��: _�TXv�B`�CEM����M3T�rC����r�_�DIAG~�RAILAC�S�bM( LO60��\6���$PSb"�� X�P`e,cPR�PS��J]�ǂC�Q� 	YC�FUN�>RINE�����r�脤10�S_����lP��pzT�d�zTCBL���&�B�A;�7q>�7�D�A!0�|�B�;�LD@�t0�Q��W!������TI��ĕ&A�$CE_RIAu�V�AF�`P��,R@��T2��C�.b��AOI�p�FDF_aL���2��LM�C}Fr�HRDYO�!z@RG��H��!��|��C�MULSE3�t�c�g3�$J�:�J�2�7�;FAN_�ALM��¢WRNʥHARD��n�	Pq�2¡�q�%Y_.@�&AU�@R�t~0TO_SBR:�/�c 7�p�S��O�M/PINFe@,qb�ܚ�m�REG��NV��z�6DU N�DF9Lu�$M���p�tĦ,`�ѨصC�M�PNFAqxcON�@q� ��@|@v�����$��$Y�$&"!+ �o� ��#EG��?#t0O�ARQ \5�2��[�h��%AXE�Y'ROBV*RED&V&WR@@1_��83CSY0��0��S���WRI@@b��`ST�� W#10�0Eq ��k�e3�_ B�fAt!֤�DFPOTO}�9��R@ARYV#X�0��Fd�� FI� �#�$LINK2�GkTHw��T_��fAj�6f2��XY�Z���7��OFF�n@w��ғ�\�BT ݂��CA� ���FIEp�?�l4݂n$_J���2���Q�0�:�8f2� (��Nၢ��CZ�%DUt�ri�9��TURŠ!X˓��f�]�X��tPn�FL��@uc\�������30f2|A +1���K{ M�$\5�3�a���e���g�ORQ:�c!���a��� O�����P���ca!�����OVE��*�M ]��#���)���/����s��wa��p��AN �az�����+���   .b�������L)�LL��c!ER�!�	��!E@@P���A8��	�5�d׃��f��AXCC���F`�ay� �e��	���	e0�
�� �
���
���
��
���
1��C��	C��	 C�C�C�,C�< C�LC�\C�l�}oDEBU�c$�`��i�-!�B��AB��ȁQ�1��VvP�b 
H"c+�p%�a|'r� |'e1|'��|'��|'�� |'�|'��������y�.��LAB�n��`��SGROopn��_PB_C�qԢ3��4�%6Y1o�U5"�a6AND+�``a�Ղ"��7 _Q��в8E��8bp��NTՠ7C�0VELI��1���6?�SERVE�0>��� $��A�q!"@POuB@R��)AY�$��ASS  ���PA�N�N� E@VE�RSIT�NG.[@0�aAImp�p�NO`@AAVMՠK� 2 �E� 0  �#5WA�O�H�O�M �L	P])_�N��@�_T_;VYU \x]�_Q�_�_�_�T�@BS��:� 1�nI� < �_o0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟����� �2��R@MA�Xo��5��c  dG�INP�b�F�PRE_EXEs�!����E�kL��A�@�IOCNV��t� �^�PǦ��s��W�SwIO_̠ 1�KP@ �?Q*��\'��@?�5���J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~�������  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o�o0mG�LARMRECOV ���Y����LMDG ���8�LM?_IF �c� 5��o�o!z�oD�Vhz�}, 
 ��/r;�����!�$�E�,�i��(������ÏՏ@�NGTOL  ��� 	 A   ���G�PPINFoO �k �f�P�b�t���Y�   �r����wb��ߟɟ� ���9�#�]�G�m���ġ�ݏ��ѯ���� �+�=�O�a�s�������jPPLICAT�ION ?�������Handling�Tool � �
V9.30P/�04���
88g340���F0 ��202�����7DF3������None��F{RA�� 6=����_ACTIVE�=b  ȳ�  ~��UTOMOD����u���CHGAoPONL�� ��OUPLED 1�i� B�F�X��j߼�CUREQ �1	�k  Tt�
t�t�	����̰���xbtҤ׵��H��E���HTTHKY�� yb�߹�����C�U�g� ������������� 	��-�?�Q�c����� ������������ );M_���� ����%7 I[����� ���/!/3/E/W/ �/{/�/�/�/�/�/�/ �/??/?A?S?�?w? �?�?�?�?�?�?�?O O+O=OOO�OsO�O�O �O�O�O�O�O__'_ 9_K_�_o_�_�_�_�_ �_�_�_�_o#o5oGo �oko}o�o�o�o�o�o �o�o1C�g�y����܆�TO�������DO_CL�EAN���I�NMw  �� t��������͏ߏz�DS�PDRYRP���H	I��s�@��K�]�o� ��������ɟ۟���8�#���MAX��0��q��!�A�X0�@�=�|@���PLUGG0и1�=���PRC�B�q�u�:�,���Ox����SEGF	�K����q���K�]��o�����˯��LAP (�;��������/� A�S�e�wωϛϭϿ�>�TOTALc�����USENU(��5� ���҆�RGDISPMMC�eh�C�S�@@��5�O&�H��1�_�STRING 1�
�
�M���S��
��_I�TEM1��  n �ͼ���������(� :�L�^�p������������ ��I�/O SIGNA�L��Tryout Mode���InpR�Sim�ulated���Outd�OV�ERR%� = 1�00��In c�yclX���Prog Aborn����N�Statu�s��	Heart�beat��MH� Faul����Aler��%�%7�I[m��� ,���,��߸ *<N`r�� �����//&/88/J/�WOR��� �!�\/�/�/�/�/�/ ??(?:?L?^?p?�?��?�?�?�?�?�? NPO����&@�+OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_p{_�_�_!BDEV)N �P=O�_�_oo'o9o Ko]ooo�o�o�o�o�o��o�o�o#5GPALT�nq�/H �������� &�8�J�\�n�������p��ȏڏ\GRIF� �����:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~� ���R���*���ޯ� ��&�8�J�\�n��� ������ȿڿ����<"Ϥ�PREGr~[� ί4ςϔϦϸ����� �� ��$�6�H�Z�l��~ߐߢߴ���(��$�ARG_� D ?�	���	���  	�$(�	[�]���(�>���SBN_CONFIG7�	�\�[�u�V�C�II_SAVE � (�~�q���TC�ELLSETUP� 	�%  O�ME_IO(�(�%?MOV_H������REP��'���U�TOBACK���	�x�FRA:\H� 2�H�~��'`��H�{��� ��w� �24/06/05� 11:02:20H�?�H�����'l���Gn�����HƄ\� ,>P�t�� ����k//(/ :/L/^/��/�/�/�/p�/�/�/Ġ�  g��_J�_\ATBCKCTL.TM��-???Q?c?u?<�IN�Iqp��n��G�MESSAG���1~�|�;ODE_D����n��8O�P�?D��PAUS:@ !��	� ,,		�?�	�>OLG2OlOVO xOzO�O�O�O�O�O�O� _
_D_._@_z_���D@TSK  �!M{��?G�UPDT��0�7d�P�6XW?ZD_ENB�4j��VSTA�5	��U���XIS\�UNT �2	�{�}�� �	 o� M7v ���š�0b��N�H�V`��ovo�o�n�:v��Ġhu��Ġ��o�o�o�o03f�MET��2�V��� PUa?Z -?���>�߿4��R�?W0+?�^l�}7GB��7jt�6&ff�3`N7@Ĝ�7AUU9}SCRDCFG 1	�;]� ���{����)�;�M�t�H�Q��������� ӏ���^����?�Q� c�u����� �:���J�GR=`�P�?ؓ0N5A���	J�Ֆ�_ED�01�y� 
 �%-0EDT-Ɵ�V�z�Ġ��e@�K�I�Hʅ?�=��B���  ���2�[�8��=w䙦��Ưدn����3������ d���Kϒ���:�ȿ�4������)ά�@�^�p�ߔ��5O� �Ϝ���)�x���*�<���`��6��h�� )�D������,��7��W�4�{�)��{� ����j����8��'� K��*���G����6���9����*ͨZl��CR�"���X� r�$6�Zؐ%�?NO_DEL�֒�GE_UNUSE��ԔIGALLO�W 1�  � (*SYS�TEM*s	$SERV_GR;ܗ @REG�%$8�#|� NUM�*�#��-PMUC u�LAYOp|?PMPAL�05�CYC10$.7>8!0%>]3ULS�v?0�%92A�#Ls?�4�BOXORI�%C�UR_�0�-PM�CNV6�01�0M>�0T4DLI��P�?�)	*PRO�GRA�$PG�_MI%>OOa@AL(/EnOXEa@B�O�.�$FLUI_RESU=7�O�/�O�D#MR�.� ��b ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[6"�LAL_OUT ��+����WD_�ABOR>0g/�sI�TR_RTN  ���pNONgSTO��t p(�CE_RIA_ILd �u0���FCFG ��0��9�_PA�@G�P 1C��U�������Ϗ��C�� ����pC��Ce �(�@C8�e@�H��CX�U`�h�p�x�U�������R�d�v����?���HE ONFI�P���G_P�01C� �1#�� ��� �2�D�V�h����KPAUS�11͕0� Bj���͕ ��ܯ¯����6�H� .�l�R�|�����ƿؿ辿��r�M�pNFOw 1͕S� � 	��O�� �=��/HiB9�����{���H�bB/H�l�B������
B��>�3����}pz��������C���F���������=�	Y=��J�O=��C���pCOLLEWCT_=�+��rR���EN/@�u���n��NDE�����s#�1234?567890[��`�!S�Y�k��
 %�}�)���߱�߷� �����T��1�C� ��g�y��������� ,���	��t�?�Q�c� ���������������L5֯!2��� �9�IO  D����v�����TRr�2!�� �	
-���"�<���_MkORz#w� ��� �<����/�%/P+�m�{$�,��I?�����x#+�K�$(+���R=�%�ϱ/��!�"C4  A�&:�+�=�A{ C�z  B� $�B��"�  @�"��+�+�:dڍ? <#�
!5<�P!99?#3�!I=�&�-�?U3z'�ݑ/Qd��!T_DEFzA ��+%J�?�$� N�US<A��0��4KEY_TBL  ���6��	
��� !"#$%&�'()*+,-.�/d�:;<=>?�@ABC�0GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~�����������������������������������������������������������������������������A��͓���������������������������������耇�������������������s��p�0LCK�<8��0�0STA��$�_AUTO_DOr��&^SIND�<M^��R_T1h_ZW�T2�_���_�T{RL�0LETE�w��Z_SCREE�N ͚k�csc�U�MM�ENU 1(�{ <o}�?|o�%[o�o �oi�o�o�o�o&�o 5nEW�{� ����"���X� /�A���e�w���֏�� ������B��+�Q� ��a�s���������͟ ߟ�>��'�t�K�]� ���������ɯۯ(� ���^�5�G�m���}� ��ܿ��ſ����!� Z�1�Cϐ�g�y��ϝ� ���������D��-��z�Q�;c_MANU3AL�_�QDBcj�f4YDBG_ER�RL�0)Jk�C ���'�9��ѿNUMLIMc��1�%T0DBPXW�ORK 1*Jk���������SD�BTB_�Q +����#4�$oD�B_AWAY����GCP �"=�S15�_ALU�M_3�B��Y�Pe� ��_��W 1,�h 
��`���������_M�P�ISJPB�@� 	OoNTIMg��$��)�
�5��M?OTNEND�?���RECORD 1�2Jk ����#G�O����+B�� �!�)P�t ����Si�a /�:/L/^/p//�/ /�/'/�/�/ ??�/ 6?�/Z?�/~?�?�?�? #?�?G?�?k? O2ODO VO�?zO�?�OO�O�O �O�OgO_�O_�Od_ v_�_�_	_�_�_�_�_ c_o*o<o�_`oKo�_ �oo�o�o�ouo�o �o8�o\n�- �%�I��"�4� �X��|������ď�֏E�3�TOLER7ENC@�Bȉ�N��L����CSS_�CNSTCY 2�3w����ُ��� A�O�a�s��������� џߟ���'�9�K��a�o������DEV�ICE 24,� ����
��.� @�R�d�v���������HNDGD 5�,� �Cz����L/S 26ͭ��� .�@�R�d�vψϮ���PARAM 7���p�՚�
��SL?AVE 8ͽ��_CFG 9�����dMC:\��L%04d.CSV�χ�cA߆�v��A n�CHv�߱����΁߶������������������JCP���އ����_CRC_OUT� :ͭ��_N�OCOD��;��~��SGN <��#M�0�5-JUN-24? 11:46q����03q�� X�Xl����������M��Þ��j������V�ERSION ���V4.2�.10��EFLO�GIC 1=,� 	��Ё�����c�PROG_E�NBtն��ULS�4 Զc�_AC�CLIM5���Ö��WRST�JNTT~�c�M�O���ш�1INI�T >,��� �/OPT�� ?�	nG
 	�R575�Û 74*�	6�7�5W��1�2����]�~TO  ���D�^�VU DEXd�('�\PATHw A��A\J�����HCP_CLNTID ?A��� 뒃����IAG_GRP� 2C� �v� 	 @�K�@G�?����?l��>��X!*E �p/,�m!���/�.?�b�?v��"i�^?�Vm?Sݘ)�f403 6�78901234q5�"@D � F �s��@nȴ@�i�#@d�/@�_�w@Z~�@�U/@O�@I��@D(�*,	0'�@�n�pn�I1��A���q�B�4,ڠ$�'�
�21.0-@)�hs@$��@ �bN@��@�0��@�D@+j
A?S?e4�j
y0j	�>R��@�N@I�@�D�@>�y@�9��@42@.v��@(��@"��\�?�?�?�?O�8L��@Gl�@B�J@<z�@6�00�`@*&@$��@�@��LO^OpO�O�O�8=�q@0�F@�|�@33@��R@-?����?��`?�+�O�O�O_ _�2\�R�@�-@�&�@�@*0��!?�?� �d_v_�_�_�_�7 8m`oroPo�o�o2o|o �o�o�o &�o�o n�^��@�r E!1�15A�AMQ�P�.��� !�YR ���?�z�0�`-5A�FH�4�N����L4R�X�`-@w�p�p��Q�x�1-r�����@�`]0�Ahf'=H�9=�Ƨ�=�^5=�Ȯ���>��`-=�,ԏ�],�� �'�Ca0�<(�U�� 4�D"Q ���)A@&�?h%�Z��}h��� ��l���֟p�����0�B��y>��y�d��R=����=��zt�`-��G���G�`-p�p�aa`�Ť@q��"@�>b,�uBʂ `�B�B��B%�`-(�/��	'��V�fb�V����\fu!e1��c+���B��BW�B{0A�W�@���/ݿ'�<���#31=��4�Cw31>
��kд��r�4��|��C�!����B��W��B#�M�8�q�$��ϒ�) ��3�����R�6��\���X����%���"�[�j#�����8�?��Y'�����\?����}_߭�"!CT_C�ONFIG D||���eg��"!STBF_TTS
����8���E:�m�MAU ��~��MSW_CF���E/+  a0(�OCoVIEW�F_�k!��/�������� ��� ��4�F�X�j� |�������������� ��0BTfx� �+���� �>Pbt��' ����//(/� L/^/p/�/�/�/5/�/��/�/ ??$?��RCX�G�u,�!�/2>\? �?�?�?�?�?�?�?��SBL_FAUL�T HO:t�AG�PMSK�*G��TDIAG I���3�������UD1: 6789012345�B��{A��25P���O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�F�wF29=�
�O+o��TORECP`OrJ
�D ro�G3k�O�o�o�o�o �o,>Pbt ������_oo��u�UMP_OP�TION!�#N0�T�RX��'IQ�PM�E �D�Y_TEM�P  È�3�B���������U�NI=�奁L�YN_BRK J��~u�EDITOR6��<�~��_H`ENT� 1KO9  �,&IRVIS�:�?��&SU�MIR <��&?PICK ;���c&�?ʟ����� ��ܟ� �(�O�6�s� Z�������ͯ���� �'��K�2�D���h� ������ۿ¿���#�@5��Y�@�}Ϗ����EMGDI_ST�A��c᥁�NC_INFO 1L_���������������ì�1M_� ���9�,��
�d ��ߥ߷��������� �#�5�G�Y�k�}�� ������������^� $�6�H�Z�h���h��� ������������ 0BTfx��� ����p��'9 K]w������ ���/#/5/G/Y/ k/}/�/�/�/�/�/�/ �/?1?C?U?oy? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O �O�O�O�O�O?�O)_ ;_M_g?]_�_�_�_�_ �_�_�_oo%o7oIo [omoo�o�o�o�o�o �o__!3E�oq_ {������� ��/�A�S�e�w��� ������я��o� +�=�O�is������� ��͟ߟ���'�9� K�]�o���������ɯ ۯ���#�5�G�a� k�}�������ſ׿� ����1�C�U�g�y� �ϝϯ���������	� �-�?�Y�K�u߇ߙ� �߽���������)� ;�M�_�q����� ���������%�7�Q� c�m������������ ����!3EWi {�������� /A[�ew� ������// +/=/O/a/s/�/�/�/ �/�/G�??'?9? S]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�/ �O__1_K?U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�O�o) C_9_q���� �����%�7�I� [�m��������Ǐ�o �o���!�׏MW�i� {�������ß՟��� ��/�A�S�e�w��� ������ُ����� +�E�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� ������#�=�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �5�'�Q�c�u����� ����������) ;M_q���� ����-�?�I [m����� ��/!/3/E/W/i/ {/�/�/�/���/�/ ??7A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O #?�/�O�O__/?9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�O�o�o �o'_1CUgy �������	� �-�?�Q�c�u����� ���o������ ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������Ϗٯ �����)�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϵ�ǯ�������!� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy ��������� -?Qcu�� �����//)/ ;/M/_/q/�/�/��/ �/�/�/	%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�/�/�O�O�O�O ?_/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�O�O �o�o�o�o_'9 K]o����� ����#�5�G�Y� k�}����o��ŏ׏� ��1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ�����)� ;�M�_�q��������� ˿ݿ���%�7�I��[�m�ϙ� �$E�NETMODE �1N����  ��������˨�RROR�_PROG %µ�%���(���TA�BLE  ����g�yߋߙ���SE�V_NUM ��?  ��������_AUTO_ENB  �Ž���w_NO�� O�������  *�*����������+�,�>�P���FLsTR����HIS���������_ALM �1P�� ���죠+Q�������"�4�F�U�_����  ��������TCP_VER �!��!�V�$E�XTLOG_RE�Q�������SI�Z����STK	�����TOL � ��Dz���{A ��_BWDk�`@ p�l��UDIZw Q��px�ħ�qSTEP������ OP_DO�%��FDR_GR�P 1R��v�d �	��#��n&����c?���$,MT�� ��$ ����WizdBk?H�B��<z� �����//</�'/`/�A*HkAoFa>��j/���
 E�� 8��!��@R�/����/T/�/�/?�A�@� <0@�33@%�E0I3=@@1d?�?�?�?F@ �5�!�!�1�>�L��FZ!D�`��D�� BT���@���{=?� y O�?6���+B���5�Zf5�ES;A{=����E��^* ��X���w���m�.�FEATU�RE S��l ���Hand�lingTool� �E��Eng�lish Dictionary�G�4D St�@ar�d�F�EAnalo�g I/O�G�Gg�le Shift��Outo Sof�tware Up�dateYmat�ic Backu�p�IHQgroun?d Edit�@�G�Camera�@F��OCnrRndI�mMS�\ommon� calib U�IS�VnfQ�PMo�nitor�[tr~�@Reliab	P��HDHCP�Y�Za�ta Acqui�s�S�Yiagno�sDQ�Akocum�ent View�e�R�Wual C�heck Saf�ety�Q�FhanGced�V�J�esc`�FrwP�Gxt. oDIO �PfiGd�gend�`Err��PLFb�m�gs�ir��@�` [ �JFCT�N Menu|`v|�S-wTP Inp�facCu�EGig�EU~gu_Pp Ma�sk Exc�`g��gHTSpProx�y Svdd�vig�h-Spe�`Sk�i�T�u?`�`mmuwnicCPons�x�ur:ppo�AVrc�onnect 2��ncrUpstr�u�B
�3�eZat`J�Fe�DKAREL �Cmd. L�pu�a�xj�Run-T�i�`Env`�pe�l +GPsEPS/�W�GLicens�evccl�`Book�(System)��JMACROs,~�r/OffseP��H�`-P
o�MR��P�REnMechStop�qt#�+b�i�b[_�x�`�@EP��od
Pwitc�h��3�:a.���O�ptmş3��pfi�lcl2�g��ul�ti-T�piS�IP?CM fun=�;��o(dwb4�[�Regei�r�p>�ri\`�FK����@Num �SelW����` Adju�p��֡Z�tatu����^j�E�RDM Robo}t�@scove�A�;�ea,��`Fre�q Anly�wRemU��an�G;�G�Servo�`���H?SNPX b��^;SNSpCli[a��RLibr�C޿�@Q f�𰪶oɀt:p�ssag4��D�� 0"S��K��/IT}7şMILIB`�:�P� Firm+RJ�P�:sAcc`Ph[TPsTXo8�eln��}�;��A�K�orq}u
Pimula�Q4}Q��u��Pa��J��_P�Q��&�pev.�7�#Prit`��U�SB port ��PiP�`a\`��R� EVNTzߌ�n?except�`|��i��մh�mVC�Qr�r�r[�V'`���4��SѰSC��K�gSGE`�V�UI�K?Web Pl������p�dZavZDT Appl�t�J�֯��GridK�play�G�LT
)�R��.�Jc�:a �x��0�3Q200i(t��Glarm Caouse/z�ed�H�Ascii�qբL�oadc`��Upl���^yc	P����u��`.vRA?й`��D�Z�inAÞ��HNR�TL�ϬCOn�@e Hel�X?�U>�؍���T�tr�kRO_S Eth��t?��$�vz����2D��PkgGUpg�@ V"��3D Tri-t_a>A��Def#�6>Ba�de^���X�[ImĐF��[��nsp#�6��64MB DRA9Mo%#FRO./tPgell�L�]sh_!Dk/}'c�z%(PpA��,ty	Ps��	b��ݐ.k{��a�R�Mmaiu`Ի�mF����Pq+�lu��z�Sp��R�OzL� Sup��������0�`�pcro�F��W􏾿�O1ouest�rtsaF�|�L�O�z����K,Pl Bu�i,�n��APLCd,OvEV�E��CGeN�OCRG�OV�DG���O�DLS�OV�BU�_V�K��+_Y�TAOUVB__qW��nZi�_TCB�_�V{_�W0{��W�eoTC�O�Wp_�W��coTEHxo`�f�O�gm�oTE_�BUVF�_�g�_UVG�_ 1w1w[oUVHsUV�IA��v�UVLN��UMW�w?o�wC_UVN�UVP�e�;UVRUVS�������UVWߏ�S�U�VGF�)�P2�OE�� E�3�E��_D�D��E�!F#oE��D�R���7TUT��01�)�y23�)�TBGGk��S�rain/�UI�ې�HMI���pCon��b����f��
"iFÌ
&KAR3EL.�ݯTP_���5��"��+�X�O� a������������߿ ���'�T�K�]ϊ� �ϓϥϷ�������� �#�P�G�Y߆�}ߏ� �߳���������� L�C�U��y���� �������	��H�?� Q�~�u����������� ��D;Mz q������
 @7Ivm �����/�/ </3/E/r/i/{/�/�/ �/�/�/?�/?8?/? A?n?e?w?�?�?�?�? �?�?�?O4O+O=OjO aOsO�O�O�O�O�O�O �O_0_'_9_f_]_o_ �_�_�_�_�_�_�_�_ ,o#o5oboYoko}o�o �o�o�o�o�o�o( 1^Ugy��� ����$��-�Z� Q�c�u���������� �� ��)�V�M�_� q����������ݟ� ��%�R�I�[�m�� �������ٯ��� !�N�E�W�i�{����� ��޿տ����J� A�S�e�wϤϛϭ��� �������F�=�O� a�sߠߗߩ������� ���B�9�K�]�o� ������������� �>�5�G�Y�k����� ����������: 1CUg���� �� �	6-? Qc������ ��/2/)/;/M/_/ �/�/�/�/�/�/�/�/ ?.?%?7?I?[?�?? �?�?�?�?�?�?�?*O !O3OEOWO�O{O�O�O �O�O�O�O�O&__/_ A_S_�_w_�_�_�_�_ �_�_�_"oo+o=oOo |oso�o�o�o�o�o�o �o'9Kxo �������� �#�5�G�t�k�}��� ������׏���� 1�C�p�g�y������� ܟӟ��	��-�?� l�c�u�������دϯ ����)�;�h�_� q�������Կ˿ݿ
π��%�7�d�[ς��  H55�2rØ�21��R7�8��50��J61�4��ATUP��5�45��6��VCA�M��CRI��UI�F��28��NREv��52��R63���SCH��DOCV�R�CSU��869z��0��EIOC.��4��R69��ES�ET����J7��R{68��MASK�ůPRXY�7��OCO��3�ȝƺ���m3��J6��53u��H'�LCH��OP�LG��0�MHCuR��Sp�MCS���0��55��MDS�W���OP�MP�R�B�5�0��PCM�R0 �����z�5�51��511�0n��PRS��69���FRD��FREQn��MCN��93���SNBA:�(�SH�LB��M��BЭ�2���HTC��TMI�L��u�TPA��T7PTX��EL��z��u�8�ǲ���J95n!�TUT�95��wUEV��UEC��wUFR��VCC��O��VIP��CS�C!CSG-�g�I��WEB��HTTf��R68�CCG�{IG�IPGS�RC��DG�H7]5��R66Y7��R/�2�R?��%�q4��b��R64�ƷNVD��R6|�R�84�\��Y86f5�90Q��J9(�91)�7 ���!��D0�Fk(CLI����CMS�֚ �ƷSTY�TO�7vt�NN��ORS��J��_�OL�(E�ND��L�S�(F;VR��V3D��wPBV!APL��wAPV�CCG�ƷCCRq�CD�C�DL5CSBi�C�SK��CTCT!B�9��0�(C���0�8C�TC��0u7�TC�7TC��CT1EQ�J@�7TE]�J@V�TF�8F�(G�8)G�I5HH5HI���@\5H,CTM�(M)HUM�8N5HP�HP�8YR�8�(TS�8WIYn5VGFaWP2��P2��vPmX�7VP�DmXF�VP�GVPR6VT���P���VTB�7Vh�IHb��V>�H�'VK�V�y�@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O�O,O>OPObOtO�C�  H55��T|A�A�U�CR78��L50�IJ614΢IATU	d�D54u5�L6�IVCAyTn�CCRI![UI�Tv�E28"ZNRE�J�52ZR63�KS{CH�IDOCV�Z�C�U�D869�K0N�JEIO!dhU4�J�R69ZESET��K[J7[R68ށZMASK�IPR�XYB\7�JOCOBl3�L�J`�L3qj[J6�L53�ZH�l�LCHQjOPLGz�K0�jMHCRRj]S{MCS�L0!k{55�JMDSWr{v�kOP�kMPR�jt~P�l0�JPCMAZ�R0�{`�Jp�k5�1[51�0ZP�RSk69qjFR�D1ZFREQ�JM�CN�J93�JSN�BAr[�kSHLB���MЋ~Pa|2�JH{TC�JTMIL�L��ZTPA�ZTPT�X�EL��p�[8��K�@�ZJ95QZT�UT�k95qjUE�VjUECQjUF]R1ZVCC�O1zwVIP!�CSCQ��CSGaZ�PI�IW�EB�JHTT�JR�6p\�CGp�IG�P�IPGS��RCv!�DG�kH75ZWR66�7 kR�E2�jR�l�P�4qj����JR64�ZNV�DjR6 {R84�����>`�86�k9�0���[J9�l91��A�7P[>`QZD0:p�F_�CLI�| [�CMS�Z���JST�Y!�TOq�7�\N]NqjORS1zJ���BjO�OL��END�JL �S��FVR��ZV3D!�@[PB�VQ�APL�ZAP�V�jCCG�JCC�RzCD �CDL���CSB�ZCSKv�zCT@�CTB1�Q�>���Cъn�1�C�A�TCAZn���TCv�TCjCTE�Z�����TE�Z��1�TUFQ�F��G1�G1�
��H��I��~���`�WCTM��M��M!�UN��P��P1�RQ얠�TSQ�W1��V�GFQP2�P2p��n ap�VPDa�FAZVP��VPR�A�VT�K� �JVT�B��V�[IH�VXΠ����VK!�Vp� �Hx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO��C�@STD~�DLANG�D �I�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ����'�9�K�RBT�FOPTNb�t������� ��Ο�����(�:�L��EDPN�Dp��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾���������*�}HH�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ������1�C�U��g�y�99~��$�FEAT_ADD ?	��������  	 }Ⱦ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j��|�������DEMO� S��   }��ݏ��� %�R�I�[�������� ���ٟ���!�N� E�W���{�������ޯ կ����J�A�S� ��w�������ڿѿ� ���F�=�O�|�s� �ϟϩ��������� �B�9�K�x�o߁ߛ� ������������>� 5�G�t�k�}����� ��������:�1�C� p�g�y�����������  ��	6-?lc u������� 2);h_q� ������/./ %/7/d/[/m/�/�/�/ �/�/�/�/�/*?!?3? `?W?i?�?�?�?�?�? �?�?�?&OO/O\OSO eOO�O�O�O�O�O�O �O"__+_X_O_a_{_ �_�_�_�_�_�_�_o o'oToKo]owo�o�o �o�o�o�o�o# PGYs}��� ������L�C� U�o�y�������܏ӏ ��	��H�?�Q�k� u�������؟ϟ�� ��D�;�M�g�q��� ����ԯ˯ݯ
��� @�7�I�c�m������� пǿٿ����<�3� E�_�iϖύϟ����� ������8�/�A�[� eߒ߉ߛ��߿����� ���4�+�=�W�a�� ������������� 0�'�9�S�]������� ������������,# 5OY�}��� ����(1K U�y����� ��$//-/G/Q/~/ u/�/�/�/�/�/�/�/  ??)?C?M?z?q?�? �?�?�?�?�?�?OO %O?OIOvOmOO�O�O �O�O�O�O__!_;_ E_r_i_{_�_�_�_�_ �_�_ooo7oAono eowo�o�o�o�o�o�o 3=jas �������� �/�9�f�]�o����� ��ҏɏۏ����+� 5�b�Y�k�������Ο şן����'�1�^� U�g�������ʯ��ӯ  ���	�#�-�Z�Q�c� ������ƿ��Ͽ��� ��)�V�M�_όσ� ���Ϲ��������� %�R�I�[߈�ߑ߾� �����������!�N� E�W��{������ ��������J�A�S� ��w������������� ��F=O|s ������� B9Kxo�� �����//>/ 5/G/t/k/}/�/�/�/ �/�/�/??:?1?C? p?g?y?�?�?�?�?�? �?�?	O6O-O?OlOcO uO�O�O�O�O�O�O�O _2_)_;_h___q_�_ �_�_�_�_�_�_o.o %o7odo[omo�o�o�o �o�o�o�o�o*!3 `Wi����� ���&��/�\�S� e�������ȏ��я� ��"��+�X�O�a��� ����ğ��͟��� �'�T�K�]������� ����ɯ����#� P�G�Y���}������� ſ߿����L�C� Uς�yϋϸϯ����� ���	��H�?�Q�~� u߇ߴ߽߫������ ��D�;�M�z�q�� ��������
��� @�7�I�v�m������ ��������<3�Eri{���  ��� );M_q�� �����//%/ 7/I/[/m//�/�/�/ �/�/�/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o�o#5 GYk}���� �����1�C�U� g�y���������ӏ� ��	��-�?�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o�������|��ɉ  ʈ ρ���	��-�?�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������΁Ӏƈ����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ ASew������	�$FEAT_�DEMOIN  ����� ��INDEX���� ILECO�MP T���7�-�SETUP2 �U7A� � N l*_AP2BCK 1V7?  �)��"�%��� :� ���*/�N/�[/ �//�/7/�/�/m/? �/&?8?�/\?�/�?�? !?�?E?�?i?�?O�? 4O�?XOjO�?�OO�O �OSO�OwO__�OB_ �Of_�Os_�_+_�_O_ �_�_�_o�_>oPo�_ too�o�o9o�o]o�o �o�o(�oL�op� �5��k �� $�6��Z��~���� ��C�؏g������2� ��V�h�������� Q��u�
����@�ϟ d�󟈯��)���M�� �������<�N�ݯr�����%���̿FzP�~ 2�*.cVRӿϋ�* ��Fψ�L�p�Z��PC�xϡϋ�FR6:D����\��π�T �'߶��Q�� ��w�Y�*.F
Ϩߊ�	�Ö���d��߈�STM�.�»��"Y���}��HJ���?��[�m����GIF�6�A�"��������JPG����A��0c�u�
��JS=⋰��+��%
J�avaScripti��CSZ�@���k %Cas�cading S�tyle She�ets�_�
AR�GNAME.DT�D�\0�P�`q`DISP*gJD�������
TPEI?NS.XML$/��:\8/�XCus�tom Tool�bary/�PAS�SWORD�}��FRS:\�/{/ �%Passwo�rd Config�/X�F?�/??|?�� �?/?�?�?e?�?�?O 0O�?TO�?xOOO�O =O�OaO�O_�O,_�O P_b_�O�__�_�_K_ �_o_o�_�_:o�_^o �_Wo�o#o�oGo�o�o }o�o6H�ol�o �1�U�y�  ��D��h�z�	��� -�ԏc�������� ��R��v��o���;� П_������*���N� `�����7�I�ޯ m������8�ǯ\�� ����!���E�ڿ�{� ϟ�4�ÿտj����� χ���S���w��� ��B���f�x�ߜ�+� ��O�a��߅���� P���t����9��� ]������(���L��� ������5�����k�  ��$6��Z��~ ��C�gy �2�+h�� ��Q�u
//� @/�d/�/�/)/�/ M/�/�/�/?�/<?N? �/r??�?�?7?�?[? �??�?&O�?JO�?CO �OO�O3O�O�OiO�O �O"_4_�OX_�O|__�_�_�V�$FIL�E_DGBCK �1V���P��� < ��)
SUMMA�RY.DG�_h\�MD:�_0otP�Diag Sum�mary1o>Z
C?ONSLOG&o	o�ato�oCaCon�sole log��o=[	TPACC�N�o%�o4?e�TP Accou�ntin�o>ZF�R6:IPKDM�P.ZIPhlX
���@ePpException�n{`�MEMCHECK�*�oo@��aMe�mory Dat�aA��V-l�)+�RIPE�o�+����O�%�� Packet L�o��TL�$��r��S�TAT������H�� %܂Sta�tusI���	FTAP����/���K��a�mment TB�D͟�� >I)ETHERNE�य़�q�P�CaEt�hern��`fi�gura�DT��DCSVRF�������үY��� verify allկޖSM.���DIFFʯ��¯W�փ�diffY���q��CHG01N�5�G�`ܿ[�o���-?��2ҿ��˿`�k���¡�3V�=�O��� �v�ߚ�VTR�NDIAG.LS������h�S�(� �Opex�� Han�osticu���)VDEV,�DATi�F�X�j�\��Vis��Dev�ice�ߟ�IMG@,ү����n�Ճ��Imag��U�P��ES��I�FORS:\����Da�Updates OList��>Z\��FLEXEVEN�F�M�_�x�[�;� ?UIF Ev����R,�s�)
P�SRBWLD.C	M��h\������`�PS_ROBOW�EL�:GIG���Wb�{N�Gi�gE����RN�?� )lHADO�Wv[mQ�S�hadow Ch�angej�w�b��RCMERR�����Q�KC�FG Error�
�tail) M�A��CMSGLIB~ew/���d��ic��7�)�ZDGf/���/M�ZD� a�d,/��NOT�I��i/{/?O�N?otificy��/���AGJ_g?n_�? �_�?�?D_�?t?	OO �??O�?cOuOO�O(O �O�O^O�O�O_�O$_ M_�Oq_ _�_�_6_�_ Z_�_o�_%o�_Io[o �_oo�o2o�o�oho �o�o!3�oW�o{ ��@��v� �/��<�e����� ����N��r����� =�̏a�s����&��� J�ȟ񟀟���9�K� ڟo�������4�ɯX� �����#���G�֯T� }����0�ſ׿f��� ���1���U��yϋ� ϯ�>���b���	ߘ� -߼�Q�c��χ�߫� ��L���p����;� ��_���l��$��H� ����~����7�I��� m������2���V��� z���!��E��i{ 
�.��d�� /�S�w� �<�`�/�+/ �O/a/��//�/�/ J/�/n/?�/?9?�/ ]?�/�?�?"?�?F?�? �?|?O�?5OGO�?kO��?�OO�O�O�C�$�FILE_FRS�PRT  ����@�����HMDONLY� 1V�E�@ �
 �)MD:�_VDAEXTP.ZZZ�O}OT_c[�6%NO �Back fil�e ._�DS�6P ZO�_D_�_�O�_oTO 3o�_Woio�_�oo�o �oRo�ovo�oA �oe�or�*�N �����=�O�� s������8�͏\�� ����'���K�ڏo��� ���4�ɟ۟j������#�5��DVISBC�KX�AS*.V�D6����FR:�\O�ION\DA�TA\k����Vision VD�R��������*� �N�ݯ_������7� ̿޿m�ϑ�&ϵ�ǿ \�뿀ϒ�M϶�E��� i���ߟ�4���X�j� �ώ�߲�A�S���w� ����B���f���w� ��+���O����������>�����t��JLU�I_CONFIG7 W�Eb�� $ ]��C������� $6T$ |xf�hz�� ��V��+ �<as���@ ���//'/�K/ ]/o/�/�/�/</�/�/ �/�/?#?�/G?Y?k? }?�?�?8?�?�?�?�? OO�?COUOgOyO�O �O4O�O�O�O�O	__ �O?_Q_c_u_�__�_ �_�_�_�_o�_)o;o Mo_oqo�oo�o�o�o �o�o�o%7I[ m����� ��!�3�E�W�i�{� �����ÏՏ����� �/�A�S�e�w���� ����џ�z����+� =�O�a����������� ͯ߯v���'�9�K� ]�����������ɿۿ r����#�5�G�Y�� }Ϗϡϳ�����n��� ��1�C�U���yߋ� �߯�����j���	�� -�?���P�u���� ��T�������)�;� ��_�q���������P� ����%7��[ m���L�� �!3�Wi{ ���D���/�///�  x�;/H#�$FLUI�_DATA X����x!��j$RESU_LT 2Yx%�  �T��W/ �/�/�/�/??)?;? M?_?q?�?�?��/�? �?�?�?OO)O;OMO@_OqO�O�O�O�M?�0��x%�O�K��_"_4_F_X_ j_|_�_�_�_�_�_�_ �3�Oo$o6oHoZolo ~o�o�o�o�o�o�o�{ �Ow�O0�OW i{������ ���/�A�Re�w� ��������я���� �+�=��o^� ��D ����͟ߟ���'� 9�K�]�o�����R��� ɯۯ����#�5�G� Y�k�}���N���r�Կ ������1�C�U�g� yϋϝϯ������Ϥ� 	��-�?�Q�c�u߇� �߽߫����ߠ��Ŀ &�8���_�q���� ����������%�7� ��[�m���������� ������!3��<� �`�L���� �/ASew �H������/ /+/=/O/a/s/�/D �h�/�/�??'? 9?K?]?o?�?�?�?�? �?�?��?O#O5OGO YOkO}O�O�O�O�O�O �/�/�/�/._�/U_g_ y_�_�_�_�_�_�_�_ 	oo-o�?Qocouo�o �o�o�o�o�o�o );�O__�B_� ������%�7� I�[�m��>o����Ǐ ُ����!�3�E�W� i�{���L^pҟ� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿�� �$� �K�]�oρϓϥϷ� ���������#�5�F� Y�k�}ߏߡ߳����� ������1��R�� v�8ϝ���������� 	��-�?�Q�c�u��� F߫��������� );M_q�B� f����%7 I[m���� ����/!/3/E/W/ i/{/�/�/�/�/�/� �/�?,?�S?e?w? �?�?�?�?�?�?�?O O+O�OOaOsO�O�O �O�O�O�O�O__'_ �/0?
?T_~_@?�_�_ �_�_�_�_o#o5oGo Yoko}o<O�o�o�o�o �o�o1CUg y8_�_\_���_� 	��-�?�Q�c�u��� ������Ϗ�o��� )�;�M�_�q������� ��˟����"�� I�[�m��������ǯ ٯ����!���E�W� i�{�������ÿտ� ����/�� ��t� 6��ϭϿ�������� �+�=�O�a�s�2��� �߻���������'� 9�K�]�o��@�R�d� ��������#�5�G� Y�k�}����������� ����1CUg y�������� ����?Qcu� ������// )/:M/_/q/�/�/�/ �/�/�/�/??%?� F?j?,�?�?�?�? �?�?�?O!O3OEOWO iO{O:/�O�O�O�O�O �O__/_A_S_e_w_ 6?�_Z?�_~?�_�_o o+o=oOoaoso�o�o �o�o�o�O�o' 9K]o���� ��_��_� ��oG� Y�k�}�������ŏ׏ ������oC�U�g� y���������ӟ��� 	���$��H�r�4� ������ϯ���� )�;�M�_�q�0����� ��˿ݿ���%�7� I�[�m�,�v�P����� �������!�3�E�W� i�{ߍߟ߱��߂��� ����/�A�S�e�w� �����~ϐϢϴ� ���=�O�a�s����� ������������ 9K]o���� ����#���� �h*������ ��//1/C/U/g/ &�/�/�/�/�/�/�/ 	??-???Q?c?u?4 FX�?|�?�?OO )O;OMO_OqO�O�O�O �Ox/�O�O__%_7_ I_[_m__�_�_�_�_ �?�_�?o�?3oEoWo io{o�o�o�o�o�o�o �o.oASew �������� ��_:��_^� o���� ����͏ߏ���'� 9�K�]�o�.������ ɟ۟����#�5�G� Y�k�*���N���r�t� �����1�C�U�g� y�������������� 	��-�?�Q�c�uχ� �ϫϽ�|��Ϡ��� ؿ;�M�_�q߃ߕߧ� ����������ҿ7� I�[�m������� ������������<� f�(ߍ����������� ��/ASe$� ������� +=Oa �j�D� ��z���//'/ 9/K/]/o/�/�/�/�/ v�/�/�/?#?5?G? Y?k?}?�?�?�?r� ��
O�1OCOUOgO yO�O�O�O�O�O�O�O 	_�/-_?_Q_c_u_�_ �_�_�_�_�_�_oo �?�?�?\oO�o�o�o �o�o�o�o%7 I[_���� ����!�3�E�W� i�(o:oLo��poՏ� ����/�A�S�e�w� ������l������ �+�=�O�a�s����� ����z�ܯ�� �'� 9�K�]�o��������� ɿۿ����"�5�G� Y�k�}Ϗϡϳ����� �����̯.��R�� yߋߝ߯��������� 	��-�?�Q�c�"χ� ������������ )�;�M�_�߀�Bߤ� f�h�����%7 I[m���t� ���!3EW i{���p���� �/�//A/S/e/w/ �/�/�/�/�/�/�/? �+?=?O?a?s?�?�? �?�?�?�?�?O�/ �0OZO/�O�O�O�O �O�O�O�O_#_5_G_ Y_?}_�_�_�_�_�_ �_�_oo1oCoUoO ^O8O�o�onO�o�o�o 	-?Qcu� ��j_����� )�;�M�_�q������� foxo�o�o���o%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ���ʏ܏�P��w� ��������ѿ���� �+�=�O��sυϗ� �ϻ���������'� 9�K�]��.�@���d� ���������#�5�G� Y�k�}���`ϲ��� ������1�C�U�g� y�������n������� ��-?Qcu� ������ );M_q��� ����/��"/�� F/m//�/�/�/�/ �/�/�/?!?3?E?W? {?�?�?�?�?�?�? �?OO/OAOSO/tO 6/�OZ/\O�O�O�O_ _+_=_O_a_s_�_�_ �_h?�_�_�_oo'o 9oKo]ooo�o�o�odO �o�O�o�o�_#5G Yk}����� ���_�1�C�U�g� y���������ӏ��� �o �o$�N�u��� ������ϟ���� )�;�M��q������� ��˯ݯ���%�7� I��R�,�v���b�ǿ ٿ����!�3�E�W� i�{ύϟ�^������� ����/�A�S�e�w� �ߛ�Z�l�~����ߴ� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������������D �k}����� ��1C�g y������� 	//-/?/Q/"4 �/X�/�/�/�/?? )?;?M?_?q?�?�?T �?�?�?�?OO%O7O IO[OmOO�O�Ob/�O �/�O�/_!_3_E_W_ i_{_�_�_�_�_�_�_ �_
_o/oAoSoeowo �o�o�o�o�o�o�o�O �O:�Oas�� �������'� 9�K�
oo��������� ɏۏ����#�5�G� h�*��NP�şן �����1�C�U�g� y�����\���ӯ��� 	��-�?�Q�c�u��� ��X���|�޿𿴯� )�;�M�_�qσϕϧ� �������Ϯ��%�7� I�[�m�ߑߣߵ��� ���ߪ���ο�B�� i�{���������� ����/�A� �e�w� �������������� +=��F� �j� V����' 9K]o��R�� ����/#/5/G/ Y/k/}/�/N`r� �/�??1?C?U?g? y?�?�?�?�?�?�?� 	OO-O?OQOcOuO�O �O�O�O�O�O�O�/�/ �/8_�/__q_�_�_�_ �_�_�_�_oo%o7o �?[omoo�o�o�o�o �o�o�o!3E_ _(_�L_���� ���/�A�S�e�w� ��Ho����я���� �+�=�O�a�s����� V��zܟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ 鿨�
�̟.��U�g� yϋϝϯ��������� 	��-�?���c�u߇� �߽߫��������� )�;���\�π�B�D� ����������%�7� I�[�m����Pߵ��� ������!3EW i{�L�p��� ��/ASew ��������/ /+/=/O/a/s/�/�/ �/�/�/�/���? 6?�]?o?�?�?�?�? �?�?�?�?O#O5O� YOkO}O�O�O�O�O�O �O�O__1_�/:?? ^_�_J?�_�_�_�_�_ 	oo-o?oQocouo�o FO�o�o�o�o�o );M_q�B_T_ f_x_��_��%�7� I�[�m��������Ǐ ُ�o���!�3�E�W� i�{�������ß՟� ���,��S�e�w� ��������ѯ���� �+��O�a�s����� ����Ϳ߿���'� 9���
��~�@��Ϸ� ���������#�5�G� Y�k�}�<��߳����� ������1�C�U�g� y��JϬ�n������ 	��-�?�Q�c�u��� ������������ );M_q��� ��������"�� I[m���� ���/!/3/��W/ i/{/�/�/�/�/�/�/ �/??/?�P?t? 68?�?�?�?�?�?O O+O=OOOaOsO�OD/ �O�O�O�O�O__'_ 9_K_]_o_�_@?�_d? �_�_�O�_o#o5oGo Yoko}o�o�o�o�o�o �O�o1CUg y������_�_ �_ �*��_Q�c�u��� ������Ϗ���� )��oM�_�q������� ��˟ݟ���%�� .��R�|�>�����ǯ ٯ����!�3�E�W� i�{�:�����ÿտ� ����/�A�S�e�w� 6�H�Z�l��ϐ���� �+�=�O�a�s߅ߗ� �߻��ߌ�����'� 9�K�]�o����� ����ϬϾ� ���G� Y�k�}����������� ������CUg y������� 	-�����r4� ������// )/;/M/_/q/0�/�/ �/�/�/�/??%?7? I?[?m??>�?b�? ��?�?O!O3OEOWO iO{O�O�O�O�O�O�? �O__/_A_S_e_w_ �_�_�_�_�_�?�_�? o�?=oOoaoso�o�o �o�o�o�o�o' �OK]o���� �����#��_D� oh�*o,�����ŏ׏ �����1�C�U�g� y�8������ӟ��� 	��-�?�Q�c�u�4� ��X���̯����� )�;�M�_�q������� ��˿�����%�7� I�[�m�ϑϣϵ��� ��Я������E�W� i�{ߍߟ߱������� ����ܿA�S�e�w� ������������ ���"���F�p�2ߗ� ����������' 9K]o.��� ����#5G Yk*�<�N�`���� ��//1/C/U/g/ y/�/�/�/�/��/�/ 	??-???Q?c?u?�? �?�?�?�?���O �;OMO_OqO�O�O�O �O�O�O�O__�/7_ I_[_m__�_�_�_�_ �_�_�_o!o�?�?O fo(O�o�o�o�o�o�o �o/ASe$_ v������� �+�=�O�a�s�2o�� Vo��zoߏ���'� 9�K�]�o��������� ɟڏ����#�5�G� Y�k�}�������ů�� 毨�
�̏1�C�U�g� y���������ӿ��� 	��ڟ?�Q�c�uχ� �ϫϽ��������� ֯8���\�� ߕߧ� ����������%�7� I�[�m�,ϑ����� �������!�3�E�W� i�(ߊ�L߮������� ��/ASew ����~��� +=Oas�� ��z������/�� 9/K/]/o/�/�/�/�/ �/�/�/�/?�5?G? Y?k?}?�?�?�?�?�? �?�?O�/�:OdO &/�O�O�O�O�O�O�O 	__-_?_Q_c_"?�_ �_�_�_�_�_�_oo )o;oMo_oO0OBOTO �oxO�o�o%7 I[m���t_ ����!�3�E�W� i�{�������Ï�o�o �o��o/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���ԏ ���Z���������� ɿۿ����#�5�G� Y��jϏϡϳ����� ������1�C�U�g� &���J���n������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��x���������%7 I[m���� �����3EW i{������ �/��,/��P// �/�/�/�/�/�/�/? ?+?=?O?a? �?�? �?�?�?�?�?OO'O 9OKO]O/~O@/�O�O x?�O�O�O_#_5_G_ Y_k_}_�_�_�_r?�_ �_�_oo1oCoUogo yo�o�o�onO�O�O�o �O-?Qcu� ��������_ )�;�M�_�q������� ��ˏݏ���o
�o .�X��������ǟ ٟ����!�3�E�W� �{�������ïկ� ����/�A�S��$� 6�H���l�ѿ���� �+�=�O�a�sυϗ� ��h���������'� 9�K�]�o߁ߓߥ߷� v������߾�#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	������N�u� ������ );M�^��� ����//%/7/ I/[/|/>�/b�/ �/�/�/?!?3?E?W? i?{?�?�?�?�/�?�? �?OO/OAOSOeOwO �O�O�Ol/�O�/�O�/ _+_=_O_a_s_�_�_ �_�_�_�_�_o�?'o 9oKo]ooo�o�o�o�o �o�o�o�o�O �OD _}����� ����1�C�U�o y���������ӏ��� 	��-�?�Q�r�4 ����l�ϟ���� )�;�M�_�q������� f�˯ݯ���%�7� I�[�m������b��� ��п����!�3�E�W� i�{ύϟϱ������� �ϸ��/�A�S�e�w� �ߛ߭߿������ߴ� ��ؿ"�L��s��� �����������'� 9�K�
�o��������� ��������#5G ��*�<�`��� ��1CUg y��\����� 	//-/?/Q/c/u/�/ �/�/j|��/�? )?;?M?_?q?�?�?�? �?�?�?�?�O%O7O IO[OmOO�O�O�O�O �O�O�O�/�/�/B_? i_{_�_�_�_�_�_�_ �_oo/oAo ORowo �o�o�o�o�o�o�o +=O_p2_� V_������'� 9�K�]�o�������� ɏۏ����#�5�G� Y�k�}�����`� 柨��1�C�U�g� y���������ӯ��� ���-�?�Q�c�u��� ������Ͽ�󿲟� ֟8�����qσϕϧ� ����������%�7� I��m�ߑߣߵ��� �������!�3�E�� f�(ϊ��`������� ����/�A�S�e�w� ����Z߿������� +=Oas�� V��z�����' 9K]o���� �����/#/5/G/ Y/k/}/�/�/�/�/�/ �/���?@?g? y?�?�?�?�?�?�?�? 	OO-O?O�cOuO�O �O�O�O�O�O�O__ )_;_�/??0?�_T? �_�_�_�_oo%o7o Io[omoo�oPO�o�o �o�o�o!3EW i{��^_p_�_� �_��/�A�S�e�w� ��������я㏢o� �+�=�O�a�s����� ����͟ߟ��� 6��]�o��������� ɯۯ����#�5�� F�k�}�������ſ׿ �����1�C��d��&��ϖ��$FMR�2_GRP 1Z���� ��C4  B�.O�	 O��������F@ ��E������H����L��FZ!D�`��D�� BT���@����?� � L�H���6����t���5�Zf�5�ES���A�3  �߮�BH���~��@�33@���	��H���������@�����U���<��z�<�ڔ=�7�<�
;;�*�<����8ۧ�9k'V�8��8����7ג	8(�� 4��X���������;�M���_CFG [��T��w�����|��O�NO ��/
F0�� ��L��RM_CHKTYP  ��O������w���ROM��_MsIN O���. u���X��SSB]��\�� ��[O�R{�S��TP_DEF_O/W  O��â�IRCOM ���$GENOVRD�_DO#Y��T[HR# d�d�o_ENB� � �RAVC��]DO  ��œ~,�Ģ����� ��FOU��c������ȷ��< + ^�8/�0/R/�/O�C�  D� �/"&d�/�,@���,B�����"��#)�GSMT°�dT��Q �$�$�HOSTC]�1e���P �Y��� kMCO��+{?�O�  27.0z�01�?  e�? �?
OO.O<J�?_OqO��O�O�<OOIC	anonymous�O �O�O_ _2_ z?��GXG[�?�O�_�?�_ �_�_�_oKO(o:oLo ^o�_o�O�o�o�o�o �o5_�oY_k_Ho�_ _����o�� � �2�U�o�oz��� ����	-?A� .�uR�d�v������ ��П����)�_� � N�`�r�����ݏ�� ޯ��I�&�8�J�\� ����������ȿ�m� 3��"�4�F�Xϟ��� ïկ׿�������� �0�w�T�f�xߊߜ� �����������,� sυϗ�t�ߘ��ϼ� ������߯�(�:�L� ^�����ߦ������� ��5�G�Y�k�m�?�� ~�������  2U����z�����/4]1ENT� 1f+ P!\K	/  +0� 4/#/X//|/?/�/c/ �/�/�/�/�/?�/B? ?f?)?�?M?_?�?�? �?�?O�?,O�?ObO %O�OIO�OmO�O�O�O _�O(_�OL__p_3_ |_W_�_�_�_�_�_o �_6o�_Zoo/o�oSo�owo�o�jQUICC0�o�o�o4�dA15#��d2��as�!ROU�TER���$�!?PCJOG%� ��!192.168.0.10�o~�cCAMPRTu�Q�!e�1n������RT������ !�Softwar�e Operat�or Panel���b�c��NAME� !�!RO�BO��k�S_CF�G 1e� ��Auto�-started^FTP'�� >@'�tK�]�o��� �����ɯۯ���� ��5�G�Y�k�}���՟ ���ֿ�/���0� B�T��xϊϜϮ��� �e�����,�>�P� );�ϼ���� ����(���L�^�p� ����9������� � �$�k�}ߏ�l���� �ߴ���������  2DVy���u�� ���-�?�Q�c�e R��v����� ��//*/M�`/ r/�/�/�/�/% ?9/&?mJ?\?n?�? G/=?�?�?�?�??O �?4OFOXOjO|O�/�/ �/�/�?�O/?__0_ B_T_Ox_�_�_�_�_ �Oe_�_oo,o>oPo �O�O�Oio�_�o_�o �o(�_L^p ��o�9��� �����z�_ERR �g��"�2�PDU�SIZ  �p^��`�I�>b�WR�D ?Õ�a� � guest�v����Ə؏����s�SCD_GR�OUP 3hÜ uǑ�yIFTB�w$PAB�OMPB�w B�_SHB��ED�� $CB�C�OM4�TTP_A�UTH 1iA�� <!iPen�dan����Ʒ!�KAREL:*8��.�KCC�S��e�;�VISION SET,�ï��4�گȯ��:�� #�p�G�Y�{�}�������CTRL j�A����q
��FFF9E3����dFRS:DE�FAULT!��FANUC We�b Server !����┊���ʼ����ϻ�������0�WR�_CONFIG �k1�}��!�2�IDL_CP�U_PC@��qB�ȕ`c� BHI�M�INT�9�g�GNR_IO;�p��pG�K��NPT_SIM_�DO����STA�L_SCRN�� ������TPMOD�NTOL�ף�|�R�TY��cѨַ��E�NB��9�H�OL_NK 1lA�>� k�}��������O�_MASTE��?����OSLAVE �mA��RAMCOACHE����O�O_CFG7�N�O��UO Z�K�CMT�_OP@���E���Y�CL6�i�:�_AS�G 1n&�|�
 ���� 2DV hz������\����NUMo�E��
K�IP4�F�RTRY_CN��i���O_UPDo�j��I�1 K�v�T�o�6���6�K�P_MEMBERS 2p&�� $1����S���K�RCA_A�CC 2q1� � X�_Q 	��S  t� 6y_� 6p,�p���A&6ϐ  3�Q/C% �rr,�#$BUF001 �2r1�= \`�u0  u0\o��$��$��$��$���$��$��$��$�V�#]44&4U64G4X4j4Uz4�4�4�4U�4�4�4��#�^�4�4/�4A��4Q�4c�4s�4���4��4��4��4��4ڄ4��#_u0�c�_�4�$�4<u0�]{H_�0�dhC ���p�[U�#[f�,Dv,D�,D�,D��,D�,D�,D�,D�,D��$
�$�$,J�$=�$N�#�)2�/ �#�!�!�B� �B� �B � �B� �B� �B� �B 0�B0�!1R0R #0R+0R30R;0R C0RK0RS0R[0R�c0Rk0Rs0i�=�z1t �1�! �1�R�0�R�0�R�0�R �0�R�0�R�0�R�0�R �0�R�0�R�0�R�0�R��0�R�0�!�1tp ��A�R@b@t� �Ac$@%@*A�! 2A7b;@7bC@7bK@7b S@7b[@7bc@7bk@7b s@7b{@�B�@�B�@�B��@�B�@�B�@�!�)3 �O�%�C�b�"�C�b�" �C�b�"S�b2S�q 3!S r#21S r32AS  rC2QS rS2aS rc2 qS rs2P{2P�2�S �r�2�S�r�2�S�r�2 �S�r�2�S�r�2�S�r �2�S�r�2c��Bc ��@���t"D2b8�3B Ac8�CBQc8�SBac8� cBqc8�sB�c�b�B�c��b�B�c�b�B�fU�2s1� 4��Ś�
�!<��������#$�HIS�"u1� ��A! 2024�-06-05�� i�Z�l�~���C ��� ��ǟٟ럸����G� 4�F�X�j�|������� į֯����0�B� T�f�x���������� �����,�>�P�b� tφϽ�Ͽ�������� ��(�:�L�^ߕϧ� �Ϧ߸������� �� $�6�H�ߑ�~��� ����������� �� �@�/�A�w�����������d������ Q�c�M_q��� ����&8J7 I[m���� �"/!/3/E/W/ i/{/�/�/�/���/ �/??/?A?S?e?w? �?�/�/�?�?�?�?O O+O=OOOaO�?�?nO �O�O�O�O�O__'_ 9_'�9�`B�T�f��_ �_�_�_�����_oo )o;ouO�Oqo�o�o�o �o�o�o�oJo\o no[m���� ���4F3�E�W� i�{�������ÏՏ� ���/�A�S�e�w� ������������� �+�=�O�a�s����� Ο��ͯ߯���'��9�K�]�K_A_I_�CFG 2vh[� H
Cycl�e Time���Busy��Idyl����mink�=ݱUp�����Read��gDowѸͿ �}��Count���	Num �����ȗ�N̉P%�3�PR�OG��whUrP�^ϣϵ����������ع.�SDT_ISOLC  hY�� =�n�J23�_DSP_ENB�  0�ްQ�IN�C xa݉S>�A�   ?�  =���<#�
=�>��:�o �Ѽ�`�߉Q����J�OBy��CZ�ٵ���G_�GROUP 1yv0���<��P�ә�\���?������PQ��������� �0�B�T�������G_IN_AUT�O�e�POSRE��*�KANJI_�MASK������R�ELMON zh[VωRy�2DV�hzn���}�{���lӉT���m�KCwL_L��NUM^���$KEYLOGOGING� mP�P��i�t�LANGUA_GE hU8��DEFAUgLT FVQLG���|��ݲ�Qx��а  8ްH�  ��P'0���P;�P�]ಉU;���
�(UT13:\�� �� �//+/=/O/f/s/ą/�.(!�/QVLN�_DISP }�{�ڸ����$OCT3OL'0�QDzn�9����=1GBOOK ~Wd�$౨!�!u0X��?�?�?�?��?�;Mc޳I�6	[5�X��]Oߎ��Y2_BUFF 2�0� ���P2 ٵ�Ot2��O׷�O�O __$_Q_H_Z_�_~_ �_�_�_�_�_�_oo� oMonӈADCS ��ɇҜ�LQO������o�o�o�oddIOw 2�pk ��!X��$4FX l|������ ���0�D�T�f�x����������ԏ�eER/_ITM-�dr�-� ?�Q�c�u��������� ϟ����)�;�M��_�q�����77�SE�V� a���TYP-�����!������RST�beSCRN_FL 2�}n���o������˿0ݿ��2�TP-���1=NGNAMpZԎ58`dUPS� SGIJ���i�p��_LOAD�G �%.�%SUM�IR��MAXU�ALRM���1@��i�
��v�_PRD{ļ� O3A��C� �e=/��O�u1��6�P 2�e; ؟&	쯚߅߾ߩ� ��������<��1� r�]��������� �����	�J�5�n�Y� ���������������� "F1j|_� ������	 BT7xc�� ����/,//P/ ;/t/W/i/�/�/�/�/ �/?�/(??L?/?A? �?m?�?�?�?�?�? O��?$O��DBGDEF � Չa,�<D�_LDXDISA�[�-��cMEMO_{APU�E ?.�
 RAH�O�O��O�O�O__,_��F�RQ_CFG �� �VCA G@i�sS@<�dd%/\Л_@_RPh҈ ��D*�P/�R **:�RD�_ �X�_Fo,oYoPobo �o�o�o�oO ��o�`�o'w,(�o l�dZ�~��� ����9�K�2�o��V�������ɏ��IS�C 1�.��P � O�DWO'�O`�K����Տ�_MSTR� �����SCD 1��M�|���x� ��>�)�b�M�_��� �������˯��� :�%�^�I���m����� ʿ��ǿ ��$��H� 3�l�W�|Ϣύ��ϱ� �������2��/�h� Sߌ�w߰ߛ��߿��� 
���.��R�=�v�a� ������������ �<�'�L�r�]����������������MK�UQ����Q$M�LTARMTR�:�W? 0sP@�~�?@METPU�y@������ND�SP_ADCOLx�T@�CMNT� �FN� ��FSTLI��� ���Uu�Qm|w�POSCF#=�PRPM���ST� 1��� 4R#�
���� /'�//#/e/G/ Y/�/}/�/�/�/�/? �/�/=??1?s?]1��SING_CHK�  $MODASS��=?�5�DEV 	|J	�MC:�<HSI�ZEyM��ȭ5TA�SK %|J%$�12345678�9 NO`E�7TRI�G 1��� l ?E�_�O6y�O�O6}0F�YPA6u�4�3E�M_INF 1���[`)AT?&FV0E0�OY]�)AQE0V1&�A3&B1&D2�&S0&C1S0}=H])ATZY_�_�TH�_�_hQ�Oo�XA	o1o�_Uo<oyo�o ?_�oc_u_�_�_ 
�_.eoRdo� C�����o�o� �o�o�o`�k%��� ��u��������8� J��n�!�3�E�W�ȟ {��#���"�ՏF�� j�|�c���S�e�֯�� �����0��T���x� 3�=���i�ҿ����� ��,�߯�����9� �ϼ���ϓ�߿���:�!�^��?NITO�R>G ?�;  � 	EXEC�1���2��3��4���5��q@��7��8
��9����(��� ���������� ������������2�2�2+�2�7�2C�2O�2[�2�g�2s�2�3�3��3�ҭ1R_GRP_SV 1�.[� (e1�C���?���� ��� \����?C���=8A_D���Ng�ION_D�B�0��=��  ��q TՅ��&����q ��8T�N�   #ߵ�\>�9-ud1E�/A�PL_NA_ME !?Ej ��!Defau�lt Perso�nality (�from FD)���RR2%� 1��L�XL�ypj�� dh �����#5 GYk}��������//1/�32 �\/n/�/�/�/�/�/�/�/�/�2<K/(?:? L?^?p?�?�?�?�?�?(�?�?I6?(N
OLOKP;OxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_UOgO �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �_�_ $6HZ l~��������� � H��6 H�b H\y�KA�  �M�_�KdI�1�~���t� ����2�%�H
�����8�+�.� �F� <�N�`�~�����ğA�Д����K�	`�0�*�<�N��:��oA�n�������? A�  ��� گ�����1�诀U�g�R���v���NRN$� 1�b	���@ � TҜj � @D[���?����?K �KA��6Ez  "��	4�;�	l�	� �@� 0<�� O� ���� �? � �t�A��J��K ���J˷�J� ��J�4�JR�<�������^���A�@��S�@�;fA�6A��A?1UA��X�ϸ���=�N��f������T;f���X�������*  ��  �5��>@��[��?���?+�?����#�K�'��ߣ��ߔ�������-�1ϻ���Є���(  +��������֢����	'� �� 2�I� ��  �ƥ��:��ÈV�È=����n���� �<O�� �� � � ���������x���� �  '�����@!�p@�Wa�@#�@'�@+�[C?�CP��P�K�B��CS�����@��  ��ɚ�0�0�ɹ�i�i���@K ��KD'�� �� $H3��s����� :Η  }��x?�ffя��X ����8��#1>�Aצ������^Ph��	e�^�^���>�������<2�!<�"7�<L��<�`N<D��<���,��������N��?fff�?��?& ޔ@T��"!?�`?Uȩ?X�2! ��z�!�Z��f/� �/�J���/�/�/�/ ?�/&??J?\?G?�?��O%F��o?�?k?��?W/O{)�?4O�8H�mN H[���G?� F��=OvO �OsO�O�O�O�O�O�O ___N_��o_yS;_ ���?�_O�_W_oo ,o>o�Soeo�_�o�o�o�o�o�o��{�
r©{C�o?�ocN}�f��mt�����e���}{�BHP�E�\��Z܉r��p��q*�@I��}@�n�@��@�: @l��?�٧]� ���%�n�������=�=D�ɋ�g���@��oA�&{C/?� @�U����+J8��
H���>��=3H���_�� F��6�G��E��A5F�ĮE���֏耎�fG���E��+E��EX�����>\�G�Z�E�M�F�lD�
��(��s�^� ��������ߟʟ��  �9�$�]�H���l��� ����ۯƯ���#�� G�2�k�V�h�����ſ ���Կ����C�.� g�Rϋ�vϯϚ��Ͼ� ��	���-��Q�<�u� `߅߫ߖ��ߺ����� ��;�&�8�q�\�� ������������� 7�"�[�F��j�����������(��4���������3��ϩ��#q4 ��{*<#q�0+q#VhJjb���1E�䴛| ���	�� 6�$�UP�PhwQ �_��������� ���1//A/g/R/#r$j/|/�/�/�/ �/�/�v_0??T?B<eZ?d?�?�?�?�?�?�Q)�?�?OOBO�0OfOtJ  2 7H�6#vH���C�\�#vBqqpB)��p�pA#p@�O #t�s�O__�OC_�V�O�O�_�_�_�_�_*#t^D#p#p�!�#p�F#u
  �_#o5oGoYoko}o�o �o�o�o�o�o�o����Q ��R����4�$MR_CA�BLE 2�RO �@�T~�A@� ?�ptq�B�mp��p�@B�@C��p�OM�`B��Xo��C��^��mv³@��@B��@M�O
�uv�p�M7v�EC�kg���x�@���@C�p9�t{���uZ*�vg�[����*�p��@��C���r7��BV�9'�I `��sÏ�ޏ��ȏ -��6�(�"�P�F�X� ������ڟ��ğ)��2��q�Y&��������m�ү�����*�** FsO�M �Sy�������%% �2345678901S�e� P���t�T� �� �A� ��
z��not? sent ����WZTES�TFECSALG!Rw0���Ad��Q���
(�u@�~��-rE�C�U�g�y� �9UD1:\m�aintenances.xml�����   j�DEFAULTK\~FrGRP 2�7��  pRXk  ��%1st m�echanical checkz�6��d��l�u�vEERZ�߲�������ߜ<�controllerL��e�:�wD��f�x�����MC���"�8��� ����vE�U�"�4�F�X�j���C ������#����� $6��CE�g�eA�. batt�ery:���vE	�����������Supply g�reasy1!B���8<B BIvE��v������N
cabl5��
e:/L/^/p/�/@I	�Y�/�)/@�/?"?4?F?� $�/n?=�@��? �/�?�? �?�?
OY?.O}?�?�? WO�O�O�O�O�OO�O COUOgO<_N_`_r_�_ �O;_�_	_�_-_oo &o8oJo�_no�o�_�o �_�o�o�o�o_o4 �o�oj�o���� �%�I[0�T� f�x���������!� ��E��,�>�P�b��� ��Տ珼������ �(�w�L�������џ ����ʯܯ�=��a� s���;�l�~������� �ؿ'�9�K� �2�D� V�hϷ�Ϟ���� ����
��.�}�R�d� �ψ��Ϭ߾������� C��g�y�N��r�� ����	���-�?�� c�8�J�\�n������ �����)���"4 F��j�������� ���[0� f������! �EWi/P/b/t/ �/�/��/////? ?(?:?L?�/?�?�/ q?�/�?�?�? OOa? 6OHO�?lO�?�O�O�O �O�O'O�OKO]O2_�O�V_h_z_�_�_\�B	 T�_�_�_�__o 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^��p�������  ̾LQ?�  @�A 
o����F͏p2�D�V��H*v�** *Q(V!��������Ο�����(���O_HS��+�y��� ��_���ӯ�/�A�S� ��?�Q�c���o����� �������)�s� ��_�qσ�Ϳ߿�� �������%�7�Iߓ�����J�$MR_H�IST 2�(U���� 
 \�B$� 2345678�901�߼�~�p���9�O�%�����O m���H�Z������� ����3�E���i� � ����V���z������� ��AS
w.� �d����+���SKCFMAPw  (U��U"�� � 3�CONREL  ����\dEEX_CFENB�
Z�B�FNC��JOGOVLIM�qd���EKEY���%_PANp�""ERUN��+SFSPDT�YP��DSIG�N��T1MOT���E_CE_�GRP 1�(U\���P#��/��/ "?�$?M??q?�?:? �?^?�?�?�?O�?�? 7O�?[OmOTO�OHO�O �O�O�O�O�O!__E_��O:_{_2_�_V[EQ?Z_EDIT�$V�#TCOM_CF/G 1�R��_�o"o 
�Q_AR�C_��%�T_MN_MODE�&{��Z_SPLFo��UAP_CPL��o�NOCHEC�K ?R * �o�o $ 6HZl~�������wNO_WAIT_L�'�W� NT�Q�RaU��<�_ERR�!2	�Rd� �������@�j܏��a`Oj�}�q�| 	�c�_�:��<9 � ?��?�Y�?�m,�c�PA�RAMk��R�؆*�ܟǗf��� = ��(�:�B�� d�v�R������������ЫƗ�&�8�˟�\�"ODRDSP��c�&�OFFSET_CAR�PLo���DIS����S_A�a`ARK�'�YOPEN_FILE����!%a�V=`OPTION_IO/!��M_PRG %�R%$*O�a��WmOް��'ك�В���  �im��M���	� �����	���r�RG_DSBOL  ��\U���o�RIENTT5O��C�l[�A p�U�`IM_ED�Yقr�Vv�?LCT �F��RХ�%a���dj�_P�EXi`����RAT�ig d��ԗ�UOP �{�������(��L�Z��$���2�#�L�X�L�pe� ��M������������ � �2�D�V�h�z��� ������������
�2��9K]o�� ����L�( );M_q�����XY��.C�/+/X�P/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?2/D/�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�Ov? �?�O�O__%_7_I_ [_m__�_�_�_�_�_0�_}��OƗ�*o<m ��K���]ookQo�o�g�mmK��o�o�g �g#+=[a ��`����|҄�d�	`��+���:�oJ�I�[�m��>$�A�  ���o ���؏��o���3� �0�i�T���l�p�v��O��1����� ���r�@ ���*�̐ �@D�  ߑ?���ˑ?5��5�D��  Ez���� � ;�	l��	 ��@�? 0���0� �ې� � �� �U��H�0#H��G��9G�ģG?�	{Gkf�ˇ`��o�����C�?����i�D	� DO@ D����r����  �5��>�����B������ BB�Bp�{�!5���O�㯈bo�u���`��Ӈ����x�����(  ������׶����{�	'� � ��I� � � ���y�=����7�I���� �<0�� �� � A¯���������ҏ���z�NK���  '�\���ġ �C<�C�?�,�B��A����߼�߰�@������{�00 ʉ��F�F���@5��� �����������)���`�r�T�d�5�� �:������x?��ff�o���9� !�p���� �85���>�ׇ��ʊΰ?�PI�d�F�?�?����>����Ᏽ<�2�!<"7�<�L��<`N<D��<��,w��������/��?fff?��?&����@T�?��`?Uȩ?X�)[����� ʉ�G�f��+��� ������� +=(asJ����2TV�/�H�mN H[�5�G?� F��/W/ i/T/�/x/�/�/�/�/ �/�/�//?яP?Z3? ����?��?8?�?�? OO��4OFO�?yOdO�O�O�O�O��\��B���KC�O _�OD_/]?��N_U_�_y_��ç����MD�H�AХI��_�:hT�xhPgQa@I���@n�@���@: @l���?٧]�_ ���%�n��߱���=�=�D�l�Hi��@��oA�&{C/� @�Ugo� �+J8���
H��>��=�3H��_�o �F�6�G���E�A5F�ğ�E��o�`���fG��E���+E��E�X��o�`>\�G��ZE�M�F?�lD�
��	 �_T?xc��� ������>�)� b�M���q��������� ˏ��(��L�7�I� ��m�����ʟ���ٟ ��$��H�3�l�W��� {��������կ��� 2��V�A�f���w��� ��Կ�������� R�=�v�aϚυϾϩ� ��������<�'�`�@K߄�o߁ߺ�ub(wa�4���w���<�է�3�ϩ����na4 �{��na��0+#7�I�+��jbc�u�1E����|�������������x5P��PI�X1e?r���~��������������� ��"H3nb$K] �������W?�5#e;E{i0����)�����#//G/U*  �2 H�6nfHY���v#\�nfB�AL�A�@B��P�PAn`@�O�/�/�/�/??(=~3�R?d?v?�?��?�?nd�n`�n`B1n`c&ne
 �?OO(O:OLO ^OpO�O�O�O�O�O�O��Omj�1 ��3�����4�$PAR�AM_MENU �?����  DE�FPULSE�K�	WAITTMO{UTR[RCVe_� SHELL�_WRK.$CU�R_STYLPP��\OPT�!�_P�TB�_�RC�_R_DECSN]P:�l oo+oToOoaoso�o �o�o�o�o�o�o,�'QSSREL_IOD  ��W!�;u�USE_PROG %6Z%(�<sCCRiPMrW!>S�w�_HOST !F6Z!�t��zTZ���s��q �:��{_TIMEgRMv�u�'PGDEBUG�Kp6[<sGINP_�FLMSKc���T�R����PGA�� 2��A?ыCH�����TYPE3\?0 '!W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿����WORD ?	�6[
 	PR<���MAI`��gSU�QC�TE!�����	�TP�CO�L��lɐ��Lip U�����ȵudw��TRACECTL� 1���@Q� G� '�G�U ����DT �Q���$���D� � 9�@U!9��0?��0�?���?��0?��0?��=�=�=�=�@=�1�C�U�gߙ�	��U
��������U��C��C��C��UC��C��C����TMp��������Au߇ߙ߽߫�E��UE��E��E��E�ԡE����w���� }������������ ����:�
��.�L�^� p��#�5�G�Y�k�}� ��������������Qcu��� ���Acu��� ����!�/�/�/ �/�/�/??1?C?U?-�u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o�����i?��ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_��_�_�_oo)i�$�PGTRACEL�EN  (a  ��'`��=f_UP �/���lat`Xa�m`=a_CFG7 �leVc'am`�d�d�o�g|O`�j  ��e��bDEFSPD ���l&aO`��=`H_CONFI�G �leTc U'`'`d3t�Lb &a6qP�d�aRq�'`�=`IN�`T�RL ��m�a8l�egqPEu�"w�la�d2q�f=`WLID�c��m	�y�LLB 1�"y� �SuBBpB94��f Sx+��%�Vu�o << %a?�U�t�U� l�������ď�؏
� (�� �B�p�V�x���Ú>�ڟџ��W��	�F�9�K�|��yGRoP 1��|(a�@�  �[��'aA?x�D P��DV�C2��$��7t�a���2q2p��p{�M��qF�´L�.��BO� v�V�@�R���v���'a�>'oY>a���ο��� =N�=R��W�� Tύ�xϱϜ�6�������	�/��  DzT�]�'`
D߅�4ߕ� �ߦ��������'�� K�6�H��l��������)(a
V7.10beta1�d�5pB(�A�\)A�G�����>�������A���*��ff�A�?p�AaG�����#@�L�� ��o�0�������cAp��Ʋ �Bq�d��#���²�?��񾢪ffA������
oH3r&a�����6�H2lV�zKNO?W_M  �e�f��tSV �"zIrc�s�(:��^I[�'a��sM����"{ ��	~�e���x��t�d������@�a�6!>%�:/L,���qMR����T�h�Ƶ�/�+��OADBANFW�D��sST��1 �1�li4?payloa���>?)`�u)?n?M?_? �?�?�?�?�?�?O�? OO%O7OIO[OmOO��O�O�O�O_�f72�<�4�O  �<I__��33_E_W_i_74�_�_�_�_7A5�_�_�_o76,o>oPobo77o�o�o�o78�o�o�o7+MA� �0s�gOVLD  ({���2PARNUM  ;�sS�n�SCHwy �u�
��q��#.�UP�D��u&�|�2_CMP_�zp0� �'�%��ER_C;HK�����!�������RS� �/��'_MO�/�_��pe�_RES_G0�({
\���������� ՟ȟڟ����/�"�S��F�w�j�]O�2PZ� j���O��P��دݯQ� �P����Q�+`7�V� [�Q�~`v�����Q��` ��ԿٿQ�$p����Q�V 1�5�!��@`}x�THR_INR� |q�z�%d��MASS�ϛ Z��MN����M�ON_QUEUE� �5�& ���*pdN��UفN���Ȏ�END�9�5�EcXED�5�Z�BEC�|%��OPTIO"��B��PROGRAoM %��%��R���TASK_�Iyt��OCFG ���Ϫ�� �DA�TA��)�@�q� 2 @���L��������    �����"�4�����  C�C�u���������INFO��m�������! 3EWi{��� ����/AS�������m�b���l��K_#��)����ENBzp�sa��2��G#�2��� X,		��=���6/��b%N!$0�N)N)v���_EDIT ��)�/�/�WER�FLe�z��#RGA�DJ ̓*A�  5? �5���&�Ѫ��u�?�  Bz�G" �<N! ���%:r?0�(�/#3}2�/7��+	H�l[�y�<1u?O Ae��t$�6�*�0/�2 **:�2 ��?CM�u6B1E���1;I�qa?]�[O)M�M9OKO yOoO�O�O�O�O�O�O �Og__#_Q_G_Y_�_ }_�_�_�_�_?o�_�_ )oo1o�oUogo�o�o �o�o�o�o	� -?mcu��� ���[���E�;� M�Ǐq���������3� ݏ���%���I�[� ��������ǟ��� ��w�!�3�a�W�i�� ����ͯïկO���� 9�/�A���e�w�������r�	<�F�� 4�m� X��9���3[ϼ�W������7PREF ��/:~�
�%IOR�ITY�ך&��!MPDSP���*W2M��UT��3�&ODU[CT��*��v�6OG�0_TG� ��*��HIBIT�_DO�(��TOE�NT 1ѓ+ �(!AF_IN�Ew�*�5�!t�cp5�]�!u�dL��!ic�mt�{>��XY(3�v�,��!)� 	A����� ���$�� �P�7�t�[�m����� ��������(L^*��(3�/9W2`?x���3>b��ƅ	G/L��4��8�>AQ2,  �%ГN`r��%�6�Z�������3sENHANCE �
�2A�d�Z/A%�֢���(��!�!PORT_NUMx��� D��!_C?ARTREPX���>��SKSTAw���oSLGS'������Q3^�Unothingb/??Q?�c?��0TEMP �؛�o?�'0_�a_seiban ���?���?O�?,OO PO;OtO_O�O�O�O�O �O�O�O__:_%_J_ p_[_�__�_�_�_�_  o�_�_6o!oZoEo~o io�o�o�o�o�o�o�o  D/hSe����{9VERSI�VЙ��p d?isablet"w;SAVE ٛ��	2670H7K55�x�O�!J/0Q�c�� 	����$�݋ԏ�e��,�>�P�^�	�����t��_�� 1���<�Ԑ �ѵޟ�ͷ�URGE B���޿�WF���zԄ4"��W#�=�bѹ*W�RUP_DELA�Y ��-��WR_HOT %+����I/��N�R_NORMAL���Ҭ��ЧSEMI��E���QSKIP����'͓x�������� ҿ��#��1��+�=� O��s�aϗϩϻρ� �������'�9���]� K�mߓߥ߷�}����� ���#�����Y�G�}� ���g���������|��RBTIF>����9�CVTMOU��'�%�9�DC�R���h� �С�B�4B�u >-�G:Q�%�jp����J���������<2�!<"7��<L��<`N<D��<��C����I[J� ������!�3Ey7RDIO_TYPE  Ý�;QED T_C�FG �$-U�B�H%�E�b�2�n$+ �8BȖ� �*8*/��N/9/r/ ]-/�/2��/��/�� �/�/?E?3?i?W?�? w7�/�?C��?�?�?O �?/OO?OAOSO�O�? �O�?�OkO�O_�O+_ _O_=_s_�O�_�Ok_ �_g_�_�_oo%oKo 9ooo�_�o�_woQo�o �o�o�o5#Y{o ��Q�M��� ��1��U�w|�� ]�����ӏ�������	�+�a���x�E�I�NT 2៩����G;� ��ț"x5�b(f�0 �  �=�@�1�P�R�d��� ������ί����� <�"�4�r�`������� ̿���޿��8�J� 0�n�\ϒπ϶��Ϯ� ������� �F�,�j��Xߎ�+�EFPOS�1 1�n  xf��ٻ�� ��)�5������|�g� ��;���_������� ��B���f������7� I���������,�� P��M�!�E� i����L7 p�/�S�� �/�6/�Z/l// /S/�/�/�/s/�/�/  ?�/?V?�/z??�? 9?�?�?o?�?�?OO @O�?dO�?�O#O�O�O YO�O}O_�O*_<_�O �O#_�_o_�_C_�_g_ �_�_�_&o�_Jo�_no 	o�o�o?oQo�o�o�o �o4�oX�oU� )�M�q��� ��T�?�x����7� ��[����������>� ُb�t��!�[����� ��{����(�ß%�^� �������A�ʯܯw� ��ï$��H��l�����+���ƿ_���2 1��h�z���2�� V�\�z�Ϟ�9ϛ��� o��ϓ�߷�@����� ��9ߚ߅߾�Y���}� ���<���`��߄� ��C�U�g����� &���J���n�	�k��� ?���c��������� ��	jU�)�M �q��0�T �x%7q�� ��/�>/�;/t/ /�/3/�/W/�/{/�/ �/�/:?%?^?�/�?? �?A?�?�?w? O�?$O �?HO�?�?OAO�O�O �OaO�O�O_�O_D_ �Oh__�_'_�_K_]_ o_�_
o�_.o�_Ro�_ vooso�oGo�oko�o �o�o�o�or] �1�U�y�� �8��\�����-� ?�y�ڏŏ����"��� F��C�|����;�ğ�_��ο�3 1� 뿕����_�J����� ��B�˯f�ȯ���%� ��I��m���,�f� ǿ��뿆�Ϫ�3�ο 0�i�ύ�(ϱ�L��� pςϔ���/��S��� w�ߛ�6ߘ���l��� ����=�������6� ����V���z����  �9���]������� @�R�d�������#�� G��kh�<� `����� gR�&�J�n �	/�-/�Q/�u/ /"/4/n/�/�/�/�/ ?�/;?�/8?q??�? 0?�?T?�?x?�?�?�? 7O"O[O�?OO�O>O �O�OtO�O�O!_�OE_ �O�O_>_�_�_�_^_ �_�_o�_oAo�_eo  o�o$o�oHoZolo�o �o+�oO�os p�D�h���<���4 1��� ����w����ԏo� ������.�ɏR��v� ���5�G�Y�����ߟ ���<�ן`���]��� 1���U�ޯy������ ����\�G������?� ȿc�ſ����"Ͻ�F� �j���)�c��ϯ� �σ�ߧ�0���-�f� ߊ�%߮�I���m�� ����,��P���t�� ��3����i����� ��:�������3���� ��S���w� ����6 ��Z��~�=O a��� �D� he�9�]� �
/���/d/O/ �/#/�/G/�/k/�/? �/*?�/N?�/r??? 1?k?�?�?�?�?O�? 8O�?5OnO	O�O-O�O QO�OuO�O�O�O4__ X_�O|__�_;_�_�_ q_�_�_o�_Bo(�:�5 1�E��_o;o �o�o�o�_�o%�o "[�o�>� bt��!��E�� i����(���Ï^�� �����/�ʏ܏�(� ��t���H�џl����� �+�ƟO��s���� 2�D�V����ܯ��� 9�ԯ]���Z���.��� R�ۿv����������� Y�D�}�ϡ�<���`� ���ϖ�ߺ�C���g� ��&�`��߬��߀� 	��-���*�c��߇� "��F���j�|���� )��M���q����0� ����f�������7 ������0�|�P �t���3�W �{�:L^� ��/�A/�e/ / b/�/6/�/Z/�/~/? �/�/�/ ?a?L?�? ? �?D?�?h?�?O�?'O��?KO�?oOUogd6 1�roO.OhO�O�O 
_O._�OR_�OO_�_ #_�_G_�_k_�_�_�_ �_�_No9oroo�o1o �oUo�o�o�o�o8 �o\�o	U�� �u��"���X� �|����;�ď_�q� �����	�B�ݏf�� ��%�����[���� ��,�ǟٟ�%���q� ��E�ίi�򯍯�(� ïL��p����/�A� S����ٿϭ�6�ѿ Z���Wϐ�+ϴ�O��� s��ϗϩϻ���V�A� z�ߞ�9���]߿��� ����@���d���� #�]�����}���� *���'�`������� C���g�y�����& J��n	�-�� c���4�� �-�y�M�q ���0/�T/�x/�/�/�O�D7 1� �OI/[/�/?�/7?=/ [?�/??|?�?P?�? t?�?�?!O�?�?�?O {OfO�O:O�O^O�O�O �O_�OA_�Oe_ _�_ $_6_H_�_�_�_o�_ +o�_Oo�_Lo�o o�o Do�oho�o�o�o�o�o K6o
�.�R �����5��Y� ���R�����׏r� ��������U���y� ���8���\�n����� ��?�ڟc�����"� ����X��|����)� į֯�"���n���B� ˿f�ￊ��%���I� �m�ϑ�,�>�Pϊ� ����ߪ�3���W��� Tߍ�(߱�L���p��� �ߦ߸���S�>�w�� ��6��Z������ ��=���a���� �Z� ������z���'�� $]����@�<�/�$8 1��/v ��@+dj�# �G��}/�*/ �N/��/G/�/�/ �/g/�/�/?�/?J? �/n?	?�?-?�?Q?c? u?�?O�?4O�?XO�? |OOyO�OMO�OqO�O �O_�O�O�O_x_c_ �_7_�_[_�__�_o �_>o�_bo�_�o!o3o Eoo�o�o�o(�o L�oI��A� e�����H�3� l����+���O���� �����2�͏V��� �O�����ԟo����� ����R��v���� 5���Y�k�}����� <�ׯ`���������� U�޿y�ϝ�&���ӿ �π�kϤ�?���c� �χ���"߽�F���j� ߎ�)�;�M߇����� ��0���T���Q�� %��I���m�����MASK 1�����:�H��XN�O  )�G�M�M�OTE  i�  ���_CFG ������PL_�RANG��������OWER ��� SM_D�RYPRG %��	�%��S!TA�RT �a
U?ME_PRO0B���_EXEC_�ENB  ����GSPD� � �;�TDB��RMIA_O�PTION����� ��INGVE[RS`j����I_AIRPUR�� �
w���MT_"�T ���OBOT_ISO�LCg�������^%NAME�����OB_ORD_�NUM ?��H755  ��/�/�)��PC_TIMEO�UT�� x�S2�32��1�j�� LTEAC�H PENDAN�� ����64h,����Maint�enance C�ons��3?U6"�O?��No UseC=?E?�?�?�?�?8�?��"NPOp �"���n�!CH_�L� � .��	�nA9O!UD1:��O;OR!�VAIL̄!d�����SRW  �l���GER_INTVALc���P]�I�V_DATA_G�RP 2�j����/ DPP��_ ��_�Yj��_�W�_o �_+ooOo=o_oaoso �o�o�o�o�o�o %K9o]��� ������5�#� Y�G�}�k�������׏ ŏ�����/�1�C� y�g����������ӟ ���	�?�-�c�Q��� u��������ϯ�� )��M�;�]���q����n��$SAF_D?O_PULS��o�p8A��ѱ��CAN�"�c��A SC ���`X�����
>!���!~1~5!��� �_Y�k�}Ϗ� �ϳ�B��������߬1�,H8C��2�Z�!�e�dZ�uі�	�<� @���߻ߐ���։ٝ� P����_ @��T�l��4�F�X�e�T D��e���� ����������0�B� T�f�x�������OE���������  /5;��o_4-Qp*U/E
�t��Di� ���1�
  � �0*1�)����� ���,>P bt������ �//(/:/L/^/p/ �/�/�/�/�/�/�/ ?�?$?6?H?Z?l?�1� �ߕ?�?�?�?�?�?O O%Ot?H�QOcOuO�O �O�O�O�O�O�O�A5O��0��M�D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o *<N`r�� �������? 8�J�\�n��������� ȏڏEO���"�4�F� X�j�|����O'U1_�� Ο�����(�:�L� ^�p���������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω���p���t������ ��+�=�O�a�s߅� �ߩ߻�������������G�Q����@�	12�345678f�h!B!��������,����� �������#�5�G�M� ��p������������� �� $6HZl ~��_����� 0BTfx� �������/ ,/>/P/b/t/�/�/�/ �/�/�/�/??(?:? �^?p?�?�?�?�?�? �?�? OO$O6OHOZO lO~O�OO?�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�O
o o.o@oRodovo�o�o �o�o�o�o�o* <�_`r���� �����&�8�J� \�n�����Q��ȏڏ ����"�4�F�X�j� |�������ğ֟�7���
����A�S��e���Cz  B}p��   �r��2�� }� r�
���  	Ĥ�����H� �/���0��د u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ���Z����� %�7�I�[�m�ߑߣ� �����������!�3�E�W��<�0�̡p��<����y�̡  ����_��|ССt  �������_�`<��$S�CR_GRP 1��*P3� �� �<�� k�	 _7��?� P�I�1�q�`�_�\���8x���u������C���E�V������S�LR M�ate 200i�D 567890�ΠLRM- 	?LR2D 4 9�?
12343���>�7��� � ?���.��.�S����M���		����%5��#H�?��C�.�f�u�v��}���<�����/h�+�� �h��,X�_JZE�[�Bǈ��a/�_"x$[�A���/  1@<��%[�@�� �/# ?���%["H���/��*[�F@ F�`2
?/.??R?=? b?�?s?�?�?�?{�_!��!�"�?�?�?
ODB�*O�?pO[O�OO�O �O�O�O�O_�O6_!_ Z_D�jZ����W�_k�A���_�_<��!@��O>�Aj�_}�@� 4o���5gYY���uo9�A� �V�e$���`S�u<�A �o�o�oz�axH#5.�\s
�� i{�T_���9���ECLVL  �<�����`Q�@�qL_DEFA�ULT�tJ����<��HOOTSTR��a�q�MIPOWERF��p}�#�L�WFD�O� #��rRV?ENT 1��q�q�D� L!DU�M_EIP�����j!AF_IN�E�܏9�!FT$���ҏ/�!bT�� ��{�!RPC_MAIN|��^��j�ǟ��VIS䗟������!TMP�PU
�ŉd��_�!
PMON_�PROXY`�Ȇe N���&�y���f�����!RDM_SR�V��ŉg�C�!�Ra_�ƈh2���!%
��M¯i~�ۿ�!RLSYNC�ܿ�8ʿ'�!gROS��N��4��s�!
CE(�MT'COMt�ȆkbϿ�{!	��CONS�ϲǇl���!��WOASRC�Ȇm��vW�!��USBX��ƈnFߣ�!STMx���Ċo����B� ������<�a�(���� ��*SYST�EM*wPV9.3�044 ��1/9�/2020 A� �zP���� y�~��_SPD_T[����_TRQ�   
��A�XIS�� ����� 2x ��D�ETAIL_ � l$DA�TETIME{P�$ERR��DC�I�MP_VEL �  	U�TOQ~]�ANGLES]��DISTg���G_{NAB�%$L{�vD�����REC�� , ���!��2 $MRA�� �2 d��IDXrD� ���� c`�$OVER_L�IMIT]� 	�����OCCUR���  H�C?OUNTER����FZN_CFG��� 4 $EN7ABLC�ST=�D��FLAGD�DEB�UaRv��r6GR�f�  � 
�$MIN_OVR�D{P$INT_�r���FACE��SAF�MI�XED��	�R{OB��$NE��PPD��HELL�; 5$�J� BASC�RS�R_I  $qN��1]� 0�1��12T3T4�T5T6T7T8��$ROO������T_ONLY{P�$USE_ABO�7��1ACKEN�B\��IN��T_wCHK�OP_��T �_PU�'M�_@�O.�E�PNS@4���T �MN��TPFWD_KAqR[��I�REP��OPTI��E�QU�E;)��DV"Y
$�CSTOPI_AL�EX��� �C�XT M1�)2�D�� TY�SO�� NB�DI�T�RIa�!['INI8����#NRQ06� �END4$KEYSWITCHB#�W!1�$HEX BE�ATM�#PERM'_LEZ�b!EW��7�UV#F�$W"S4D�O1�M� O
�EFPS����b�5�� %C�0��E��OV�_MS!R ET_IOCM���2�&�!���HK	� D H�1SU�B�"MP�I�PO~�$FORCA#�WARN�$�O}M*  
 @;@#FU���SU��5!SAR� �E2�F3�FQ4�A����Og L�By��<(UNLO �@��DED@�(��SNPX_AS>w 0?ADDq �s$SIZC��$VAR��M�I�P�S�@A�A? � $,)P��2	APD�BC<V��VFRIFD���S� �I�4)�F34ODBUS_AD/�A�S�Y{$' ML1D�IAxA$��MY�1�!e3h4a��S2 � L0Ps�TE
d8b�SGL>aTA@  &S WcB���P`?`��T�!pcPS3EG�"paBW� @d�SHOWxeE�BA=N�`TPOF�Qd�9h0h�!��V�C� G� L`$�PC�����`��$F�B�A���fSP� A���e�aD�`�o� �;�A0�� K}�?q�@Fw�@Fw�@�Fw�@Fw5Dy6Dy7�Dy8Dy9DyADyB�Dy�@Fw �Fw�`FwF Dx�`�Py`�jy$`T��y1�y1�y1�yU1�y1�y1�y1�y1�y1�y1���ه�Py2]y2jy2wy2��y2�y2�y2�y2��y2�y2�y2�y2��y2�y2�3Cy3�Py3]y3jy3wy3��y3�y3�y3�y3��y3�y3�y3�y3��y3�y3�4Cy4�Py4]y4jy4wy4��y4�y4�y4�y4��y4�y4�y4�y4��y4�y4�5Cy5�Py5]y5jy5wy5��y5�y5�y5�y5��y5�y5�y5�y5��y5�y5�6Cy6�Py6]y6jy6wy6��y6�y6�y6�y6��y6�y6�y6�y6��y6�y6�7Cy7�Py7]y7jy7wy7��y7�y7�y7�y7��y7�y7�y7�y7��y7�y7�'BVPz�0U�� ����I
��V�R� x $TORl�!�P  _�MO�������Q_ RE�"rn��b@]�S�C4X!(�B�_U�PM��RYSL�� � 0U�RN�T%W�e ?p�0y�
rVALAUN	 \&��Fj��ID_L33��HI���IxB$FILE1_0#���$�3)`�h�SA�� h���1�E_BLCK��#>�YaG�D_CPUW�1PW�%PY���Yd`*#R ? � PW �l�P��LA~aS���������RUN_FLG��������Z0������H* ��' ���xT2\!_LI��B  #G�_O�"d P_E3DI�)pT2� GO�I�R�xP�P�m BC20t ��5`���P�GFqT�$��#TDC��A1^ � M�P��&�TH�PnQ���R� PI@ERVAE�#*�#*a����  X ;-$ULEN�#b�#U� RA� �Bi��W_#��1U��2&�MOO��ES�P�I >������U��DE��QLACE�B�CC�C>�0_�MAP�"%�"!T#CV),J!�T<1K* j%`*r�q�%�q�J� A�eM�$�0JH"7.p��!�a�2�0�P&p�!� PJK 6VK�a1a1�a0J�a*13JJv3JJ&3AAL3@L03L0F6%aJ25} N1q,}0<+& <��L�_la�0���v�CFR `��GROU��Za�Rq�N� CnS�0REQ�UIR�PEBU��SQ�&$T�2�AR�6�P�� \�@�APPR�@CL<�
$X NNKHCLO� [IS��pI�
�YV 䂉 M� ' | �B�D_MGa�@C0p2�H�p$ �GBRK�IN�OLD�F�`RTM!OFZ�M�EJF  TPN4 3 &3 j3( s3 6;U7;ULa�<R�� B|�a�Wa�SPATH�W�Q�S�Q���S�@@@��`S�CA�WLB�AINFTUC��`CpKUMhY����  $a��0?j�P?jK?`�PAYLOA�GJ{2L��R_AN��cL���i�azi�a�E�R_F2LSHR$�aLO�dba�g!c|�g!cACRL_� epgrd2H��<��$H�B2rFLE�XNC� J� P8B��);�0��JT : as��w�tv 1���F1�q)�=�������/m�E /(/:/L/^/p/�/�/ �/D�a��'�# 4Q�s� �/�/�/�q�*T��B�X*�K��%����	5� �?'?9?K0O5X5F5`j5s?�?�?�9 	Nq�4  �� �?�?�?��0��ATV� A� E�LĀ�(�HJ@v@JE�@CTRa�Q�TN��$��7HA_ND_VB<�Nqܿ��T! $��F24�F���SW�1�C��F"� $$M �`�I��Aո�A��ص)R�A��w`�F��D ɸMA�L���JA�KAA�K+��Kp��JD�K�D�KP�PG����S�T�G���I��N�HDY��I@�F�3Ř`V �g�q�g�ayg 7�����EPCULUUU^UgU�pUyU�R�2J�#1 ˰�t�R ~���<}A��ASYM�U>�	@�V"/�l�ao_& �h`,d]䜸 6oHoZolo~cJ�l6P��j���ic�_VI����}C�V_UANf���;��aJ5 2�`�2��l6��eC�g� �m� y6P)���a?tGsKr� HR� ��$����ap[D)I�@�3O N��Nӣ% K�:�I�A:Q�c4W�B�BZ�� �Pǀ�� & �� ��ME��Џ�]��D�T��PT@�๠�P��0�4`p�|����	T��1� $DUMMY}1K$PS_T��RF��P$�n�@FLA�0YP����$GLB_Tΰ��� iqΠ��U�a' X8@�7�Q�ST��@SBR��PM21_VH�T�$SV_ER�`O�o�[sCL/[A�ŀO7��GL��E�W�1( 4�0�+$Y<�Z<�W�� ��a��A^ b���U.�) ��N����$GIe�}$� (�@����1* L�0�n�}�$Fn�E&NEA�R��N[�FH)��T�ANC[���JOG�
�,P +ˠ$JOINT�����ޡMSET�1, E �E.%Ɓ�S���p"�1-� � ]�U��?�@L?OCK_FO�`��� BGLVX�GL��(TEST_XM�N@�!EMP� H�82-� $U�p�F��2)@�<1*2h��� <1(]CE�0|
#]0 $KAR�}M	TPDRA�z4q!VEC�p�6u kIU<1+A1HE� OTOOL��3V�;RE�0IS3�u�296^QQ�ACH� @E,�1O�P��3�Q�	 SI>B  �@$RAIL_B�OXE���RO�BO4?��HOWWAR:q,A� �1ROLM�RE���4�cB�@E��PO_F��!�HTML	5��a������RH��1�Q.}.�pR�0�O�r/}"��!�@�  �OU�"0 t�85(D�.���� RPO�A�PIP6N���2B�1�c�<1�@�pCORD�ED� �P�@E XT�+P�)��OD  �1 D OB`�2�� �WzQ��zRn�4�SYSzQA�DR3���� TCH�� 2 ,��E�N��jqA�!_���T����VWVA~`3 � �0����PREV_R�Tm�$EDIT�,fVSHWR�PGK`�����Do �3�bd;�$HECAD��|`��4c�KE�� CPSP]D�fJMP�PL��2��R��4�P_q��VI0S3�Cy�N�E�04�o�TICK����MhqsQ�cH=N=5 @�P�ať�a_GP*vFkpgSTY�R�1LO/P��b&r�p6�@
'`MG�U%$a�=GS)�!$(���t� 1 �P
�*vSQ�Ut0���TER�C� <���SӤ7   S槤��t�ħ1�O� }_�IZh���PR]P0�H��a�@PU��X�g_DOM"�PXS� �K��AXIw�vCA1UR�Ń4�3@pȥV���_�0�RET���P�"�P��vpFd��wpA������9 G2K���SR��8l�pι� ݺ3��E��3��3� �3�,�y�N�y�^�y� nƋ����ɋ�ɜ�ҩ�	C���Cȝg�y��ܝ���SSC 79 h�DS8p{1f� SP. ��AT\���Y�p�b�AD�DRES�3B7`S�HIF�B21_2C�H3��QI6����TU6I� :>�BCUSTOل�!V�"I";�R�(��T<���
:
�BV�A�h�b < \EX� vpG�� `��C����܂V�Vy���TX_SCREE|R=��=�qTINA� �״��Q������> T�av<��QuR�$ƅ��R�� �3`RRO7�b �P�`���a;UE�d? ����Qr� S��QRSMp�{�UfP�p������S_���!������!�⹁C�"��� 2->ҰUE��@(�\��H�GMTz�LT����b"Q�A�BB�L_�0W� b A ��S�N�O�Z�L�E�e�2@�d�RI;GHn�BRD�ߡOCKGR� ��TgP|�ג�WIDTH C�X`��A��1�I�@EY�@aB d���@Q@Zr@D�B�ACKXq�	��h FOTQ�LAB�c�?(h I�0�"$UR8AI�n ��n }HD� C 8��Bb _{a��l�o R�@�"� H�l�Z�O�Jb D!p���Uz�r��R�"]ALUM����٠ERVQsP�ЩPL ��Ef �G�EM�3!׀mR�`LP$��E�pj�))�z��7���7��06�54�6
4�74�8��r%�C�PL ����1�!S `�D��USR�'F <En U�,���FO��PRI���m@&� TRI�PAm�UND-O�dG��p$ �}�DA|���41���p �Hg���G�G pTv@X���bOS�wR��J�N�1>I����:t�41	U�>J�����9uNOFF0�K꜠�O- 1�I P?J PGU�QP>�BZU�d�ѷSUB:r vrE/_EXE�PV�aN�WON� L� �n��WA7`��z1�ՠV_DB���U�SRT� �M0!ra!�@'�OR�0 %'RAU,�$T)�Wr�_*`�dN |5���XOWNQ �T$GSRCU����pD0<l%*�MPFIQt����ESPT����5��A���2C9%E`�GO `� ��T�n�pCOP�$��S _� �2�!�A5�CT�Ӧ�#��2L �`PB/� P�SHADOW���3P1?_UNSCA�3P3���]3DGD�1�QE�GAC�#<�uQG�۲Q (�NOX���LpPE�����VW�4qGĀ�Ro � �PVEU���2ANG���6��6��2LIM_X �%F�%FH*AL��`�7 ��0�VF���#�VCCzp�dS�2C�pRA|w�0�u\�bNFA2`Z5pE�Q G��f��RRS DE�2���STEa�3�� ܣ�!��Y4� ;�)A�sp� �1+U�PP_AFP��C�@[��@�T�# Ar�Q�s�El]Ȼq��/�C��mUDRI�0lV�1V3p�T�`�+�D��MY_UBY���M��uV��p�bia�X41
bP_f0��$bL^�BMa��$�`DEY�cEXX'Qu6QMU�`XW�M��US���� _AR������6G�PACI�D�0v!�4��b�b��b��RE���>�RS�bp�U �� G�0P����`�SSR� ppV �г�C��ъ	�"u�RTSW�`�C@б0$caF�O���A�hs�3�E%�UE�3@��� SSHKZRW����z�1+�ep)��3EA�N�y��hu� SRMwRCV�X ��UO�@M�C��	�r8�c�rREF:�� ��qB�?p���zP�@�P��r���_i  �z���{�� Pa�C��R�˰�B"SR�Y ���1��5rܣ���U$GROU����c(���C�@T
uY�2��$0ذ��e 0�V��Y�X<��٠UL�AW� �C6@��XR`O�NT�#��42���᜖����[�Lcŕcŕ���ї��AT!�q�Z �t� MD�HPHUؽA�0�SA�3CM�PU�F�0�(��_���R�D��P��sЁX�c���GF?0r�[, &��M���PUF_S�1b�`0�ROx�,�;��U��L�SbURE����b3RI�c�IN�#� �?
OKt!.It!�qG�INUbH��H��V@�=B�Q���ӥ�WW��gQ�S6Sa�yfLO@�S�1P��U���NSI�D�!0�4�x�4�>HX_PE=��Yg�Z_M-S�2WD�Ys4C2���R��RSL/\ �$"�?1M ���UaCG`GtA�P�l�r�v � ��!e��h���� į֯�N��o��~����VIA�] ���HDR��J�O��"��$Z�_UP+Q�_LCOW�վ�Z�t��27LIN�EPO�� o	�Ѿ������A��pfS��^ 5^h�PATHc  h�CACH��m�
������u10�#C9AI2T�F��TD���'$HO�_"r����St��������!�PAGE�� VPx�b�@8�_SIZ�CB�ZCP=�+S@���CsMPb��AIMG�4�	�AD���"MR1E���G�GPPH`�� 6ASYNBU=F6VRTD����|G��DLE_2D=D(ɲ	C�AUAc
�yQ�p��ECCU�h�VEM�`m�T��VIRC����������LA�c�!NFO{UNo�DIAG 	RUaXYZ��Ua�W%q�H���q T�@BbIM��u0���GRABBցY\SqpLERz`CD�b߂FS�=��50D�͑Gۑ�pfS��_� pBACKL�AS��(�R���`�  W��T�c @��R�T$R��@��a A�1�� u���Ti� �!XQ� ���eI�Jt���B9PEVE�A��PPK�`����GI�NO�!BaPQ3p�HO� �Bb � �b���H� y&S����7�"RO�3AC�CELO�MQ�%VRo�UG�� �!Bb�06& AR�3PA� �.�[�D�3REM_Bf� ��3pJMh��&rc���$SSC��lq��
���0'd ��
�S��ƹNc4��LEX�e{ T�ENAB�xBbg�CFLDR�HFI �G���H8d�s�O�P2X�f�� $��V�a�MV_PI�C�4H�P��@�P%�IF�/RZ J;D3E@H�$HH�3E��1GARE��LOOS��JCB�J'2��CON8�SPLA!N� ��"C�F+Ut/�)I��GMpa�KTUFS�PUa�E+QH��E@gG�-�4 LRH��!�< RKx��!VAN9C�3kR_O���0g (�=�L��c8#$���R_A?@�0h 4��_�^p� �n�D�Q�0i �h~p+9��n��OF	F, ��g� �� ���EA%�
��< SK���M`�VIE�`2�h �P��0�j < �:脯��������pD�@�^��CUST��Up�k $W�TIT>-�$PRl1��OPTqlq�VS)F�p�l� �p��	��bMO��m�Y2�3�$J�`؅��u�_g��`nY2�g��_����XVR���o}�`T�%���ZABC���p �r�9�
��ZD4 CwSCH�q L�` �t� �
�5�!��ӀG�GN)��rLu���p�_FUNX���� �
�ZIP��r,Y2# LV<�L₎����ZMPCF��usrU��r�!h�D�MY_LNX`Ma �T����tt �$����m�CMCM���C<�C6���-�P~�Q $Jǃ��D-�͂ނׇېㅄې��_��<�܂�U�X�l�UXEUL -��҅&��&�8�J�x8�Z�ƀFTFLʆ܇�/��Z+�u���;zF�D1��Y�D� v 8 �$R��U�AN�EI3GH�#�h?((0yv��qv0��uw �0q �c,��p$B����Psb_SHIF,T�=xRVf F���p	$E�� C��6� d�`Ұ�1r�
�����D��TR��pV:�Q���SPH� ���x ,(0ܘ�� ��$G�I��KL �?%�����  (�%SVCPRG!1F0*�5��25�:�"$�3]�b�$�4����"$�5����$�6տڿ"$�7���$�8%�*�R$�9M�R�!�0u� {�%�'���$�O���$� w���$����$�ǿB� $��j�$�ϒ�$�?� ��$�g���L���
�L� ��2�L���Z�L�߂� L�0ߪ�L�X���L��� ��L���"�L���J�L� ��r�t� ����$�� ���D�*N 9r]����� ���8#\G n�}����� �"/4//X/C/|/g/ �/�/�/�/�/�/�/? 	?B?-?f?Q?�?�?�? �?�?�?�?O�?,OO�>ObOMO�O��݀V ����MC=:�H4���D�� 2�����b_x 	���,���O	_R�O2__V_ =_O_�_s_�_�_�_�_ �_
o�_.o@o'odoKo �o�o�O�ouo�o�o�o �o<N5rY� }������&� �J��o?���7����� ȏڏ�����"�4�� X�?�|���u�����֟ ��ϟ�c�0�B�)�f� M���q��������˯ ���>�%�b�t�[� �����ο%�򿩿� (��L�3�pς�iϦ� ���ϱ��� ���$�� H�Z�A�~�տsߴ�k� �߿������2��V� h�O��s������� ��
����@���d�v� ]��������������� ��<N5rY� �����Y�& �J\C�g�� ������4// X/?/|/�/u/�/	�/ �/�/?�/0?B?)?f? M?�?�?�?�?�?�?�? �?OO>O%O7OtO{Cd �{F	bO�O�O��O�O�O�O_&[%�x&_K_RS���dQ QdUt_�Wl_�_�_�_ �_�_�Y8_o`Y�_Jo 8ono\o~o�o�o�o
o �o.o�o"F4j Xz�o�o��� ���B�0�f���� �V���R�Џ���� �>���e���.����� ����̟����X�=� |��p�^��������� ȯ�0��T�ޯH�6� l�Z���~�����ۿ� ��ƿ���D�2�h�V� ��ο���|������� ��
�@�.�dߦϋ��� T߾߬���������� <�~�c��,���� ��������D�j�;�z� �n�\����������� �@���4��Dj X�|����� �0@fT� ���z��/� ,//</b/��/�R/ �/�/�/�/?�/(?j/ O?a??:??�?�?�? �?�? OB?'Of?�?ZO HOjOlO~O�O�O�OO �O>O�O2_ _V_D_f_ h_z_�_�O�__�_
o �_.ooRo@obo�_�_ �o�_�o�o�o�o* N�ou�o>�: �����&�hM� ����n�������ڏ ȏ��@�%�d��X�F� |�j�������֟��� <�Ɵ0��T�B�x�f� ��ޟïկ�������� ,��P�>�t�����گ d�ο��޿��(�� Lώ�sϲ�<Ϧϔ��� ��������$�f�Kߊ� �~�lߢߐ��ߴ��� ,�R�#�b���V�D�z� h��������(�� ���,�R�@�v�d��� ���� ������� (N<r�����b ����$J �q�:���� ��/R7/I/ /"/ �j/�/�/�/�/�/*/ ?N/�/B?0?R?T?f? �?�?�??�?&?�?O O>O,ONOPObO�O�? �O�?�O�O�O__:_ (_J_�O�O�_�Op_�_ �_�_�_o o6ox_]o �_&o�o"o�o�o�o�o �oPo5to�ohV �z����(� L�@�.�d�R���v� ���� ��$����� <�*�`�N���Ə���� t���p�ޟ��8�&� \�����L�����Ư ȯگ���4�v�[��� $���|�����¿Ŀֿ �N�3�r���f�Tϊ� xϮϜϾ��:��J� ��>�,�b�P߆�tߪ� ����ߚ����:� (�^�L���ߩ���r� ���� ����6�$�Z� �����J��������� ����2t�Y��" �z�����: 1�
�R�v ����6�*/ /:/</N/�/r/�/� �//�/?�/&??6? 8?J?�?�/�?�/p?�? �?�?�?"OO2O�?�? O�?XO�O�O�O�O�O �O_`OE_�O_x_
_ �_�_�_�_�_�_8_o \_�_Po>otobo�o�o �o�oo�o4o�o( L:p^���o� � ��$��H�6� l������\�~�X�Ə ��� ��D���k��� 4������������ �^�C����v�d��� ����������6��Z� �N�<�r�`������� ��"��2�̿&��J� 8�n�\ϒ�Կ������ ��~���"��F�4�j� �ϑ���Z��߲����� ����B��i��2� ������������� \�A���
�t�b����� ������"����� ��:p^����� �� "$6 lZ������ �/�/ /2/h/� �/�X/�/�/�/�/
? �/?p/�/g?�/@?�? �?�?�?�?�?OH?-O l?�?`O�?pO�O�O�O �O�O O_DO�O8_&_ \_J_l_�_�_�_�O�_ _�_o�_4o"oXoFo ho�o�_�o�_~o�o�o �o0T�o{� Df@����� ,�nS�����t��� ������Ώ�F�+�j� �^�L���p������� ܟ��B�̟6�$�Z� H�~�l����
�ۯ� �����2� �V�D�z� �����j�Կf��
� ��.��Rϔ�yϸ�B� �Ϛ��Ͼ������*� l�Qߐ�߄�rߨߖ� �ߺ����D�)�h��� \�J��n�����
� ��������"�X�F� |�j������������ ��
TBx�� ���h���� P�w�@� �����/X~ O/�(/�/p/�/�/�/ �/�/0/?T/�/H?�/ X?~?l?�?�?�??�? ,?�? OODO2OTOzO hO�O�?�OO�O�O�O _
_@_._P_v_�O�_ �Of_�_�_�_�_oo <o~_couo,oNo(o�o �o�o�o�oVo;zo��a�$SERV_MAIL  �e�zp�`xOUTP�UToxz�`@dtRV 2v�`}p (qJ��dtSAVE�|~yTOP10 2�y d �o6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я������*�u�YP�asF�ZN_CFG u}s�t�q��uj�GRP 2�t�� ,B  � A���aD;� �B���  B4~�sRB21�voHELLm�u��v�p����,�%RSR,�-�?�x� cϜχ��ϫ������� ��>�)�b�M߆ߘ�~���  �z�`�����߸��� �`1��������҅2�`d��U�߶H�K 1	�  ����������� �.�)�;�M�v�q��������������ټOM�M 
�-޲FTOV_ENBot��q�um�OW_RE�G_UIMbrIM�IOFWDL x���WAITJAN録��pn�t�	TIMn����VAnp��_U�NITI�yLC�g TRYn�u�dpMON_ALI_AS ?e	�phe5����� �//'/9/�]/o/ �/�/�/P/�/�/�/�/ ?�/5?G?Y?k?}?(? �?�?�?�?�?�?OO 1OCO�?gOyO�O�O�O ZO�O�O�O	__�O?_ Q_c_u_�_2_�_�_�_ �_�_oo)o;oMo�_ qo�o�o�o�odo�o�o %�oI[m *������� !�3�E�W��{����� ��Ïn������/� ڏS�e�w���4����� џ������+�=�O� a����������ͯx� ���'�ү8�]�o� ����>���ɿۿ��� ��#�5�G�Y�k�Ϗ� �ϳ����ς����� 1���U�g�yߋߝ�H� ��������	��-�?� Q�c�u� ������ z�����)�;���_� q�������R������� ��7I[m *������ !3E�i{������$SMON�_DEFPROG &����� &*SYSTEM*�~� $JO��RECALL ?�}� ( �}�5copy fr�s:orderf�il.dat v�irt:\tem�p\=>10.1�09.3.132?:18788�}/܏/�/ }-7&*.dK/]-e/�/??�&�
xyzrate 61 �/�/�/w?�?�?�%77P?j0V? h?�?OO�#87/I(?mpbackO?�?�}O�O�O }/7Bmdb� *LO^OgO�O�
__�$3x7D:\ �OAP�O�@�O|_�_�_
� 47Ua?_Q_�El_ �_o!o4OFO�O�O{o �o�o�OMo�Oho�o 0_�_�_f_w�� �_?Q�_����?~�?19552 ���y������#tp?disc 0A�S��T�f���	���%t�pconn 0  ��ҏ�u�����,o>o �oH�����o�oӟ K��x�����/@�� P�k���� ��į֯�S��}����� }|7�cd5984 U� g���
�ϯ$��˷ ӿ�vψϚ�-�?�N��`�����(?:211 ������w߉ߛ߮%�.7�:pick.tpD?ǻf���	�� ����Ұ����x��� /߿�S�e�����-� ?�����t��������O�a���)���sumir��ľ��x ��/�S��Vh� �����w� ���Rd�// ,>��s/�/�/� �N/`/�/??(/:/ �/�/o?�?�?�/�/J? \?n?�?O�?6?�?�? �?}O�O�O�?FOXOjO�O__��7��ɟ�O4#__�_$_��>�Y_���g_�_
oo#c�$�SNPX_ASG 2���Ba��  �0��%�#ojo  �?�3fPARAM� BeLa W�	XkPmd��9mh�d�C`5`�OFT_KB_CFG  mcHe2c�OPIN_SIMW  Bk�b�);Es5`RVNO�RDY_DO  ��e�eWrQST_P_DSB~�b|�*kSR Bi � &�j��w��t�cTOP_ON_ERRd3b	��PTN Be�<��A&�RI?NG_PRM�vr�VCNT_GP �2Be�aO`x 	�������������.gVDk�RP 1v�a�`ҁBqď� .�@�R�d��������� ��П�����*�Q� N�`�r���������̯ ޯ���&�8�J�\� n���������ݿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�i�f�xߊߜ� �����������/�,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZ� ~�������  GDVhz� �����/
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�?��?�?��PRG_CoOUNT�f�<�NIENBQ�EMAC��dNO_UPD 1}�{T  
O 0R�O�O�O�O�O�O_ -_(_:_L_u_p_�_�_ �_�_�_�_o oo$o MoHoZolo�o�o�o�o �o�o�o�o% 2D mhz����� ��
��E�@�R�d� ��������ՏЏ�� ��*�<�e�`�r��� ������̟����� =�8�J�\��������� ͯȯگ���"�4� ]�X�j�|�������Ŀ �����5�0�B�L�_INFO 1��El@��	� eϩϔ��ϸ�@�9�@?k�<���>�Ϻ��/H�iB9�����{��HџbB/Hl�����? AҀ��K�� C�����
B��>��3���}pz����\����C��F���������=�	Y�=�J@YSDOEBUG&@�@�\��doI��SP_PA�SS&EB?��L_OG ���A�  \�K�b� � �kA\�UD�1:\��i���_M�PC�݆EW�i�A��� �A7�SAV ��5A����ⶉ��SV.�T�EM_TIME �1���@ 0�\�f����hD��MEMBK  �E�kA����k�}���wX|l@� @����Я��������	%
�� ��@ 
�M_q��ϧ� ����, >Pbt�����<e��//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?��SKB�G�1AV��?�?��?��7\�FI2t��+�A�>  �[�����&O3I('!��;kO�:�O�����` ��O�H0�O_#_G_C�l_~_�_�_�_\�$�_�_�o o%o7oIo[omoo�o �o�o�o�o�o�o!�3EWK?T1SV�GUNSPD�� �'���zp2MO�DE_LIM ����vt2�p�q�I���uuASK_OPTION��J�����q_DI��EN�B  0��� �B�C2_GRP 2�i5��	�B���9PC�Y@X�n|BCCFGg /��� ������`��*��Ώ ���=�(�a�L��� p�������ߟʟ�� '��K�6�[���l��� ��ɯ���د�#�+��=��p�����_� ����ܿǿ ώ� �L� ��(�N�<�r�`ϖτ� �Ϩ���������8� &�\�J߀�nߐ߶ߤ� ��������"��2�4� F�|�b�M�������� ��b�����>�,�b� t���T����������� ��L:p^ �������  6$ZHjl~ ������/ /2/ D/�h/V/x/�/�/�/ �/�/�/
?�/.??R? @?b?d?v?�?�?�?�? �?�?OO(ONO<OrO `O�O�O�O�O�O�O�O __8_�P_b_�_�_ �_"_�_�_�_�_�_"o 4oFoojoXo�o|o�o �o�o�o�o�o0 TBxf���� �����*�,�>� t�b���N_����� ���(��8�^�L��� ����t�ʟ���ܟ�  �"�$�6�l�Z���~� ����دƯ����2�  �V�D�z�h������� Կ¿�����"�@�R� d�⿈�vϘϾϬ��� �����*��N�<�r� `߂߄ߖ��ߺ����� ��8�&�H�n�\�� �������������� 4�"�X��p������� ��B�������B Tf4�x��� ����,P> tb������ �//:/(/J/L/^/ �/�/�/n��/�/ ?? $?�/H?6?X?~?l?�?��6�0�$TBCS�G_GRP 2��5� � ��1 
 ?�  �?�?�?!OO EO/OAO{OeO�O�K�2��3�<d@ ���A?�1	 HB�L�H�0�F�DB$  C��2_&X�O_�Cz&_n]AбH3�33?&ff?���EA�_�_~P �H���V�U�P3DH�_�]@��P�E0�Qe�DaD"�A9o o�_(o�oLjX�FX �e�o�o�o�o�o�o�:Wf{<x�q	�V3.00�2	�lr2dfs	*`�p�t�2�p �q�<y �p�}�  a�#�2��1J2�3��=�qd�A�CFG�  �5�1 ��0h�����h�������� �0���;�&�_�J� ��n�������ݟȟ� �%��I�4�Y��j� ����ǯ���֯��� �E�0�i�T������2 � ����οx���� 7�"�[�F��jϣϵ� ���ϔ�����!��1� W��1�?|߈?�ߎߠ� ����������B�0� R�x�f�������� �������>�,�b�P� ��t����������� ��(:�/Rd� ������  "HZl*|~� ����/ /�D/ 2/h/V/x/z/�/�/�/ �/�/
?�/.??>?d? R?�?v?�?�?�?�?�? �?�?*OONO<OrO`O �O�O�O�Ov�O�O_ �O8_&_H_J_\_�_�_ �_�_�_�_�_o�_4o "oXoFoho�o�o�olo �o�o�o�o0T Bdfx���� ����*�P�>�t� b���������̏Ώ�� ��:�(�^�p�_�� ��X�V�ܟʟ ��$� �4�6�H�~�����`� ��دƯ��� �2�D� V��z�h�������Կ ¿����
�@�.�P� R�dϚψϾϬ����� ����<�*�`�N߄� rߨߖ߸ߺ����|� �,�>���n�\�~�� ����������"�4� F��j�X���|����� ��������B0 fT�x���� ��,<>P �t������ /(//L/:/p/^/�/ �/P�/�/V�/? ? 6?$?Z?H?j?�?~?�? �?�?�?�?O�?2O O VOhOzO�OFO�O�O�O �O�O
_�O.__R_@_ v_d_�_�_�_�_�_�_ �_oo(o*o<oro`o �o�o�o�o�o�o�o 8�/�/btL ������"�� F�X�j�|�:������� ��ď����0��T� B�x�f����������� �����>�,�b�P� r����������ί� ���(�^�L���p� ����ʿܿ����� ¿H�6�l�Z�|�~ϐ� �ϴ������ ���D��2�h�Vߌ�v�  �ж� ���߶���$TBJOP_�GRP 2!~���  K?���	����#������@�� 0��  � � � � ���� @���	 ߐBL  f�C�� D����[������<�B�$\����@��?�33C�p� ��~�����f�x����*�;�2��♙�@��?� �zX���s�AЄ�Ȇ � ��S��>�������;��p�AW�?�ff@&?ff?�ff����~� �����;7�I
:v,�?L������DH$ { ��@�33�"4��>������8��a��Z�O�D"� #����ZVh9���� ��������/ =//�\/v/`/n/�/ �/�/b/�/?�/�/,?L]?��C���O���	V3.09�	�lr2d�*�0�Ѷ?�7 �E8� EJ� �E\� En@ �E�E�� E��� E�� E��� E�h E��H E�0 E�� E��0�� �E��0� E��x E�X F���2D�  D��` E�0P �E�0$�00@;��0G�0R@^p �Ek�0u��0@��0@�(�0� E���0��0�X 9��IRzAF<�E�*(�ߦO�B���CV�����O��ESTPA�RS�@������HR�PABLE 1$*���@���H�GQ *��I�G�H�H��׽��G	�H
�H��HKU���H�H8�H�A+SRDI3_��J_\_n_�_�_�UdOo&k0oBoTofoxn,RSo�� �Z9K ]o������ ���#�5�G�Y�k� }�����p��IWЉ �o�o�o�o�_�_�_�_��_�X,R��NUM [ ~���B���� �@�@,R_CFG %��L�Z��@��IMEBF_�TTQG���$P�V�ER�C����R� 1&;[ 8$�?����T� ��ۏ  <�N�`�r����� ����̯ޯ���&� 8�J�\�n���ɿ���� ��ڿ���"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� x��ߜ߮��������߀��,�>�P�R$�_ԙ��@�PMI__CHAN� �} ��DBGLV�����Q��ETHERAD ?U���@d�b�*�x<�X��ROUT�!�j!p��a�?SNMASK��>�255.���3��������3POOL�OFS_DIP�����ORQCTRL '+��c�OlT[������ � 2DVhz ����Z��/�SPE_DETA�I��1
PGL_C�ONFIG -�������/ce�ll/$CID$/grp1/�/�/�/�/�/c�W��/? ?*?<?N?�/r?�?�? �?�?�?[?�?OO&O 8OJO�?�?�O�O�O�O �O�OiO�O_"_4_F_ X_�O|_�_�_�_�_�_ e_w_oo0oBoTofoڎ}�_�o�o�o�o�o �od���m��_S ew����_�� ���+��O�a�s� ��������J�ߏ�� �'�9�ȏ]�o����� ����F�۟����#� 5�G�֟k�}������� ůT������1�C� үg�y���������ӿ b���	��-�?�Q�� uχϙϫϽ���^��π��)�;�M�_�Z ��User V�iew o)}}1�234567890�ߢߴ���������X{�O#���v�2�� ��T�f�x������}�37���� �2� D�V���w�%�4��� ��������
i�+%�5��dv�����%�6S*<@N`r��%�7 ���//&/�G/%�8��/�/�/�/�/��/9/�/2 l�Camera ��w/@?R?d?v?�?�?xbE3?�?�?�>��O�O&O8OJO\OR	   66�/?�O�O�O�O�O _�?*_<_N_�Or_�_ �_�_�_�_�/�6�� c_o*o<oNo`oro_ �o�o�oo�o�o &8�_�W���o�� �����o��&� qJ�\�n�������K �WxK=����(�:� L��p�����ߏ��ʟ ܟ� ����5�� \�n���������]�گ ���I�"�4�F�X�j� |�#��W��ȿڿ� ���"�ɯF�X�jϵ� �Ϡϲ������Ϗ��W n)�4�F�X�j�|ߎ� 5ϲ�����!����� 0�B�T����9�ߕ� ���������� �%� 7���H�m����������V*	50M� &8J\���� K�����"�� ��!0#;�{��� ��|�//hA/ S/e/w/�/�/B5�K 2/�/�/??/?A?� e?w?�?�/�?�?�?�? �?O�/���[�?SOeO wO�O�O�OT?�O�O�O @O_+_=_O_a_s_O ,Eg{
_�_�_�_�_o o�O=oOoao�_�o�o �o�o�o�o�_,EӋvo +=Oas�,o� �����'�9� K��o,E?�������� ͏ߏ��'�9����]�o���������^�  b����
�� .�@�R�d�v�������   ��ğ��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲�����������ﰬ  }
^�(  �ڐ( 	 .�d�R� ��v������������*��N�<�r�8�̪ �������� N���#5GY`� ���������� %lI[m� ������2/ !/3/zW/i/{/�/�/ �/�
/�/�/?R//? A?S?e?w?�?�/�?�? �??�?OO+O=OOO �?sO�O�O�?�O�O�O �O__\OnOK_]_o_ �O�_�_�_�_�_�_4_ o#o5o|_Yoko}o�o �o�o�_�o�o�oBo 1CUgy�o�o� ���	��-�?� Q��u��������Ϗ ����^�;�M�_� ����������˟ݟ$� 6��%�7�~�[�m�� ��������ٯ���D� !�3�E�W�i�{�¯�� ��ÿ
������/�8Aψ�h�@ c�p�Ȃϔ�c�j�N����+frh:\tp�gl\robot�s\lrm200�id��_mate=_��.xmlP��� ��0�B�T�f�xߊ��ߌ����������� ��%�7�I�[�m�� ��ߢ���������� !�3�E�W�i�{����� ����������/ ASew����� ���+=O as������ �//'/9/K/]/o/ �/��/�/�/�/�/�/ ?#?5?G?Y?k?}?�/ �?�?�?�?�?�?OO�1OCOUOgOyO�N���� jϸ�<<w �� ?��K �O�O�O�O_�O_L_ 2_d_�_h_z_�_�_�_ �_ o�_o6oo.oPo�~o����(�$T�PGL_OUTP�UT 0����;�` �e�o �o�o	-?Qc u������� ��)�;�M�_�q��e��@��`2345678901������ ̏ޏ���������1� C�U�g�y��}�����ӟ�����}�)�;� M�_�q�	������˯ ݯ�����7�I�[� m�������ǿٿ� ������3�E�W�i�{� ��%ϛ���������� ���A�S�e�w߉�!� 3߿���������� '�O�a�s���/�� �����������K� ]�o�������=����� ����#��1Yk�}��9�b $$mb{���	 �-QCug� �����/�)/ /M/?/q/c/�/�/�/�/�/�/?}�A?-? ??Q?c?u?�=@�O�?��?�J ( 	 ?�?�?OO9O'O ]OKOmOoO�O�O�O�O �O�O�O#__3_Y_G_ }_k_�_�_�_�_�_�_��_ooCo���  <<�/xo�o �`go�o�o�o�o�o�� do*<�oHrL^ ������&� 8��\�n��V���>� ��ڏ�Ə�"���
� X�j������z���֟ 4�F�����&�T�.� @���������үl��� ����>�P���X���  �r���ο����b� �:�L��pς�\ϊ� ��Ϡ��� ߚ�$�6� �"�l����Ϣߴ�N� �������� �2��6� h��T�������� D�������R�d�>� �����������|� ��$N������ 0����r 8J�6�Zl���Zb)WGL1�.XML�?��$�TPOFF_LI�M _`�0[a{�&N_SV �  �4%*P_�MON 1We�'$�0�02)S�TRTCHK �2We%&?"VT?COMPAT:(�!�)&VWVAR �3Z-�(>$ R�/ �/�0m"!�_DEFPROG� %�)%IRVISIU U?,�_DISPLAY� �./2INST_�MSK  �< �k:INUSER��/q4LCK�<�;Q?UICKMET0�?�/2SCRE@�We�"tpsc@q4�1!@&I%"7@_;I�ST�*%)RACE_CFG 4Z)��$o 	4
?���HHNL 25>:7`�A�+ 2�O�O �O_"_4_F_X_jZ�EITEM 26�K� �%$1234567890�_�U  =<�_�_�_�S  !�_k0�_Jo3�_ko�_�o �oo�o)o;o_o �o/U�o�o�o�o	 �7�	��?� ���A������Ϗ 3�ۏW�i�{���M��� q���珏����A� �e�%�7���M���� �������ů���a� 	�������#�ͯy��� ���տ9�K�]���� ��S�e�ɿq������ #���G���}�/ߡ� ��|��ϗ��ϧ���S� C�U�g߁ߋ���[� ����߷��-�?�� c��5�G���S����� ��w���)�����_� ����^��y���� �7�m-� =cu���! �E�/)/�M/� ��Y/q//�/�/A/ �/e/w/@?�/[?�/?��?�/�??+?�?�DS�B7�O�:�  uR�: �APOG9
 ]O�OjO�O(J�UD1:\�L���AR_GRP �18�[� 	 @P0�O[�O1_ _U_C_y_g^��P�_��ZsQ�O�_�_�_�U?�  o)koIo7o mo[o�oo�o�o�o�o �o�o3!WEg��	�5��	CS�CB 29K o��#�5�G�Y��k�}����<UTOR?IAL :K�O�ڏGV_CONFIG ;M�AMO��O9��OUTPU�T <I*���E���������џ �����+�=�O�a� '�v���������ѯ� ����+�=�O�a�r� ��������Ϳ߿�� �'�9�K�]�n��ϓ� �Ϸ����������#� 5�G�Y�k�|Ϗߡ߳� ����������1�C� U�g�xߋ������� ����	��-�?�Q�c� t�������������� );M_q�� ������ %7I[m~�� �����/!/3/ E/W/i/z�/�/�/�/ �/�/�/??/?A?S? e?w?�%�t��?�?�? �?�?O!O3OEOWOiO {O�O�/�O�O�O�O�O __/_A_S_e_w_�_ �O�_�_�_�_�_oo +o=oOoaoso�o�o�_ �o�o�o�o'9 K]o���o�� ����#�5�G�Y� k�}������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϴ����� �����!�3�E�W�i��{ߍߟ߂8������ߺѩ��ߞ?� 1�C�U�g�y���� ����������-�?� Q�c�u����������� �����);M_ q������� %7I[m ������� !/3/E/W/i/{/�/�/ �/�/�/�/�/?//? A?S?e?w?�?�?�?�? �?�?�?O?+O=OOO aOsO�O�O�O�O�O�O �O_O'_9_K_]_o_ �_�_�_�_�_�_�_�_ o"_5oGoYoko}o�o �o�o�o�o�o�oo 1CUgy��������	���$�TX_SCREE�N 1=��;�М}��\� n���������J�� I�����,�>�P�Ǐ ُ��������Ο��W� �{�(�:�L�^�p��� �����ʯܯ� �� $�����Z�l�~����� ��+�ؿO���� �2� D�V�Ϳz��ϰ��� ������oρ�.�@�R� d�v߈��Ϭ�#����������*��N��$�UALRM_MS�G ?8��E� F�z�������� ������.�4�e�X����|���a�SEV � o���_�E�CFG ?8��B�  u@��  A   B�t
 ��"s8� BTfx����������GRPw 2@�� 0v�	 ,Na�I_�BBL_NOTE� A��T���l"r=�$q� aDEFPRO�k�%o� (%�IRVISIONOy%����/� 8/#/\/G/�/�/}/�/��/�/XFKEYD?ATA 1B8�8Op v;�>?P?'?t?�?]:,(��?�?t(POI�NT  ]�?�> ? OOK T 	O��?NDIRECT�OO CHOIC�E�?FOTOUCHUPqOrO�O�O�O �O�O	___?_&_c_ u_\_�_�_�_�_�_�_�^9��/frh�/gui/whi�tehome.png�_<oNo`oro�o��fpoint�'o�o�o�o�o �f = elook�b�o�@Rdv�|indirec�o�����
�~choic&c�J�\�n�������`ftouchup�ʏ܏� ����dfarwrg �L�^�p�������� ß՟�������A� S�e�w�����*���ѯ �������=�O�a� s�������8�Ϳ߿� ��'϶�K�]�oρ� �ϥ�4���������� #�5�e:�a�s߅ߗ� �߻���������'� 9���]�o����� F��������#�5�G� ��k�}���������T� ����1C��U y�����b� 	-?Q�u� ����^�// )/;/M/_/��/�/�/ �/�/�/l/??%?7? I?[?�/m?�?�?�?�? �?�?z?O!O3OEOWO�iOkvK�`����O�O�M�O�O�O�F,�_(_�_L_ 3_p_�_i_�_�_�_�_ �_ o�_$o6ooZoAo ~o�owo�o�o�o�o�o �o2VhGߌ ������?
�� .�@�R�d�v������ ��Џ�􏃏�*�<� N�`�r��������̟ ޟ����&�8�J�\� n��������ȯگ� ����"�4�F�X�j�|� �����Ŀֿ���� ��0�B�T�f�xϊ�� �����������ߩ� >�P�b�t߆ߘ�'߼� ���������:�L� ^�p����}���� �� ��$�+�H�Z�l� ~�������C�������  2��Vhz� ��?���
 .@�dv��� �M��//*/</ �`/r/�/�/�/�/�/ [/�/??&?8?J?�/ n?�?�?�?�?�?W?�? �?O"O4OFOXO�?|O �O�O�O�O�OeO�O_ _0_B_T_�Ox_�_�_��_�_�_�_���[}������o@!o3moUogoAf,S �oK�o�o�o�o�o �o:L3pW�� ���� ��$�� H�/�l�~�e�����Ə ؏����� �2�D�V� e_z�������ԟ� u�
��.�@�R�d�� ��������Я�q�� �*�<�N�`�r���� ����̿޿���&� 8�J�\�n����Ϥ϶� �������ύ�"�4�F� X�j�|�ߠ߲����� ���߉��0�B�T�f� x������������ ���,�>�P�b�t��� ����������� �:L^p���� ���� $� HZl~��1� ���/ /�D/V/ h/z/�/�/�/?/�/�/ �/
??.?�/R?d?v? �?�?�?;?�?�?�?O O*O<O�?`OrO�O�O �O�OIO�O�O__&_ 8_�O\_n_�_�_�_�_ �_W_�_�_o"o4oFo �_jo|o�o�o�o�oSo �o�o0BT+ �V{�+ �����}{���v,Ï���,��P� b�I���m��������� Ǐ����:�!�^�p� W���{�����ܟ�՟ ���6�H�'l�~��� ����Ư�o���� � 2�D�V��z������� ¿Կc���
��.�@� R��vψϚϬϾ��� ��q���*�<�N�`� �τߖߨߺ�����m� ��&�8�J�\�n��� ����������{�� "�4�F�X�j������ ������������0 BTfx��� ����,>P bt�]����� �/(/:/L/^/p/ �/�/#/�/�/�/�/ ? ?�/6?H?Z?l?~?�? ?�?�?�?�?�?O O �?DOVOhOzO�O�O-O �O�O�O�O
__�O@_ R_d_v_�_�_�_;_�_ �_�_oo*o�_No`o ro�o�o�o7o�o�o�o &8�o\n� ���E���� "�4��X�j�|�����h��ď�Ƌ���������5�G�!�,3�x�+� ������ҟ����ݟ� ,��P�7�t���m��� ��ί�ǯ��(�� L�^�E���i������ ܿ� ��$�6�E�Z� l�~ϐϢϴ���U��� ��� �2�D���h�z� �ߞ߰���Q�����
� �.�@�R���v��� �����_�����*� <�N���r��������� ����m�&8J \�������� i�"4FXj �������w //0/B/T/f/��/ �/�/�/�/�/�/Ϳ? ,?>?P?b?t?{/�?�? �?�?�?�?O�?(O:O LO^OpO�OO�O�O�O �O�O _�O$_6_H_Z_ l_~_�__�_�_�_�_ �_o�_2oDoVohozo �oo�o�o�o�o�o
 �o@Rdv�� )������� <�N�`�r�������7� ̏ޏ����&���J� \�n�������3�ȟڟ@����"�4�06���0����_�q���[�������, ��诛���0�B�)� f�M������������ ��ݿ��>�P�7�t� [Ϙ�ϼ��ϵ����� �(�?L�^�p߂ߔ� �ߵ������� ��$� 6���Z�l�~���� C�������� �2��� V�h�z���������Q� ����
.@��d v����M�� *<N�r� ����[�// &/8/J/�n/�/�/�/ �/�/�/i/�/?"?4? F?X?�/|?�?�?�?�? �?e?�?OO0OBOTO fO=ߊO�O�O�O�O�O �?__,_>_P_b_t_ _�_�_�_�_�_�_�_ o(o:oLo^opo�_�o �o�o�o�o�o �o$ 6HZl~�� ����� �2�D� V�h�z������ԏ ���
���.�@�R�d� v��������П��� ����<�N�`�r��� ��%���̯ޯ��� ��8�J�\�n��������{@���{@���Ͽ��˿�'��,�X��|�c� �ϲϙ��Ͻ������ 0��T�f�Mߊ�q߮� �ߧ��������,�>� %�b�I���wO���� ������%�:�L�^� p�������5�������  $��HZl~ ��1����  2�Vhz�� �?���
//./ �R/d/v/�/�/�/�/ M/�/�/??*?<?�/ `?r?�?�?�?�?I?�? �?OO&O8OJO�?nO �O�O�O�O�OWO�O�O _"_4_F_�Oj_|_�_ �_�_�_�_���_oo 0oBoTo[_xo�o�o�o �o�o�oso,> Pb�o����� �o��(�:�L�^� p��������ʏ܏� }��$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v�������� п���ϕ�*�<�N� `�rτ�ϨϺ�����������P��>�P���?�Q� c�;߅ߗ�q�,���� {������"�	�F�-� j�|�c�������� �����0��T�;�x� _������������� �_,>Pbt��� ������ :L^p��#� ��� //�6/H/ Z/l/~/�/�/1/�/�/ �/�/? ?�/D?V?h? z?�?�?-?�?�?�?�? 
OO.O�?ROdOvO�O �O�O;O�O�O�O__ *_�ON_`_r_�_�_�_ �_I_�_�_oo&o8o �_\ono�o�o�o�oEo �o�o�o"4F j|�����o� ���0�B�T��x� ��������ҏa���� �,�>�P�ߏt����� ����Ο��o���(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z�l���������ƿؿ �y�� �2�D�V�h� ���Ϟϰ��������� ���.�@�R�d�v�� �߬߾������߃��*�<�N�`�r��[p����[p���������������,��8���\�C����� y������������� 4F-jQ��� ����B )fxW���� ���/,/>/P/b/ t/�//�/�/�/�/�/ ?�/(?:?L?^?p?�? ?�?�?�?�?�? OO �?6OHOZOlO~O�OO �O�O�O�O�O_�O2_ D_V_h_z_�_�_-_�_ �_�_�_
oo�_@oRo dovo�o�o)o�o�o�o �o*�oN`r ���7���� �&��J�\�n����� �����ڏ����"� 4�;�X�j�|������� ğS������0�B� џf�x���������O� �����,�>�P�߯ t���������ο]�� ��(�:�L�ۿpς� �Ϧϸ�����k� �� $�6�H�Z���~ߐߢ� ������g���� �2� D�V�h��ߌ����� ����u�
��.�@�R� d������������������$UI_IN�USER  ������  ����_�MENHIST �1C � ( " ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,14�����9)n�621�*�<N` l,290������	'v7//A/S/�e/�-�edi�t�IRVISION/�/�/�/�/ ��7?I?[?m?p?�48,2r?�?�?�?�?���?O-O?OQOcOuO��	Ai	O �O�O�O�O�O _O$_ 6_H_Z_l_~__�_�_ �_�_�_�_�_�_2oDo Vohozo�oo�o�o�o �o�o
�o.@Rd v�)���� ���<�N�`�r��� ���O�Ȍޏ���� &�)�J�\�n������� 3�ȟڟ����"�4� ßX�j�|�������A� ֯�����0���T� f�x���������O�� ����,�>�Ϳb�t� �ϘϪϼϧ������ �(�:�L�O�p߂ߔ� �߸���Y��� ��$� 6�H�Z���~���� ����g���� �2�D� V���z����������� ��u�
.@Rd ���������� ��*<N`ru ������� &/8/J/\/n/�//�/ �/�/�/�/�/�/"?4? F?X?j?|???�?�? �?�?�?O�?0OBOTO fOxO�OO�O�O�O�O��O_���$UI�_PANEDAT�A 1E����>Q  	��}c/frh�/cgtp/fl�exdev.st�m?_width�=0&_heig�ht=10nP_Pi�ce=TP&_l�ines=3nPc�olumns=4�nPfonvP4&_�page=dou�b_P1_�)p�rim�_�_  }��_oo1oCoUogo )io�oto�o�o�o�o �o�o/A(eL���������   ���RdQ_c_u^�2�_�_�V2��Wdual]����_���� Ώ�����(��L� ^�E���i�������ܟ ß ��$�6��Z��~�@S������į֯ ���M����B�T�f� x��������ҿ���� ݿ�,��P�7�t�[� �Ϫϑ��ϵ�����s ~�	�A�S�e�w߉� ���Ͽ�2������� +�=��a�s�Z��~� ������������9� K�2�o�V������*� ������#5��Y ��}�����> ��1UgN �r�����	/ //?/����u/�/�/ �/�/�/"/�/?x)? ;?M?_?q?�?�/�?�? �?�?�?O�?%O7OO [OBOOfO�O�O�O�O L/^/�O!_3_E_W_i_ {_�O�_?�_�_�_�_ oo�_AoSo:owo^o �o�o�o�o�o�o�o +O6s��O
_ ������h9� �_]�o���������� ɏ�ԏ���5�G�.� k�R�������ş��� ������y�)�b� t���������)P�� T�Я��1�C�U�g� ί��r��������̿ 	��-�?�&�c�Jχ���πϽ�M��s�{�$�UI_POSTY�PE  �u� 	 ��� ���QUICKM_EN  ����#���RESTOR�E 1F�u  ���BV��ߧӕ�V�m�� �� ��$�6���Z�l� ~���E��������� ����-�?���z��� ������e�����
 .@��dv��� W����O*< N`����� o�//&/8/�� W/i/��/�/�/�/�/ �/�/"?4?F?X?j?? �?�?�?�?�?�/�?�? Oy?BOTOfOxO�O-O �O�O�O�O�O_�O,_�>_P_b_t_.�SCR�E>�?C��u1sc��u2��T3�T4�T5�T6ʯT7�T8�Q�STAT��� Rӧu�ʏUSER�P�_�Tk�s�SBd3Bd4Bd5*Bd6Bd7Bd8Ba���NDO_CFG �G��9�8���PD��Q,i�N�one1�#`_IN_FO 1H�u�`P�0%z_�oM��o  DV9z�o �����
����@�'��aOFFSEOT K���aM� S��_������Ǐ� ���*�!�3�}�7��� {�������ß����@�U�S�W�E�z�
j��V�a�aWORK L�mX���ۯ��O�"`UFRAM�E  ���f�aR�TOL_ABRT8>��cV�ENB_�P�?GRP 1M��O�Cz  A��� ���a��ſ׿�����1�R�=�U��an�?MSK  ���a�n�N;�%�i�%x'���p�_EVN^�b���f�Ƅb2No��
 h�aUE�V^�!td:\�event_usger\��"�C7'�d|�PF���SP ��%�spotwe{ldW�!C6��]�o߱P��!��6��� )���j�����\�� <�N���r������ 3���W���J����� ��n�������/�� ��e��FX��|���
��WŠ2O-i��8�Yk G��}��� �/�2/D//h/z/ U/�/�/�/�/�/�/
?�?�/-?R?d?�$V�ARS_CONFuI�`Po� FPS{�k<CCRG�bCSo����?TU]D8� BHA�pG��1C�A��GA?�)@���=��ͶCAA �3MR��2�Yo�c�P	��`ڢ%1: S�C130EF2 Q*�O�@T�T����j��5P�a+AA�@CC��> ��H�O!�_(_U_zAP_}_�E/�A�0�i_�_�2 B����Q�2�Ta_�_ A_o�_Bo-ofoQo�o uo�o�oo�o�o�o�o�,�_Pb�5TCC��3Z��/A�y/�;D�w0GF|0�[o���02345678901��r��qA�1������Eq�5B�P�B�pFL@�AA:�o=L �RtEj��Aڡ�Bg�3HEA�Q�D��p b��?����"�4�/� M�S�e�w��������� я����B�=�O� u�s�������ү͟ߟ ��,�'��b�]�� ��������ɯۯ���<��tMODE�ȏ4� �tRSLT 3\�<C%"�� ���o����<��sp���|�C�tSELEC���;��qD�IA_W�O1]�5R�� �,		��Q���y�G�P ����;�=�RTSYN'CSE(Ѻ9��1���WINURL ?��s@��������,�>�P�r5ISI?ONTMOU(�u���� �h�s^Sۣ�SۥP�q FR:\j�\DATA\V� �� MC���LOG��   7UD1��EX���1�' B@ ����Gab�riel_Faria���?�c�,@7F�� n6  �������2 �-ƌ�>A  � CE�4������TRAIN�;B���d��pCE�� '#`�=��ԍ�:VB_�{ (q	 UyU_q��� ����%7\Ib�STAW�`�y@�B�@�����$�\�e�_GE�sa�{;�  �
W��0|8"'HOMIN�p_bSۮ�U ؠ�(ƱƱKAC�w���%�JMPERR 2=c�{
  Q��� �/r��3�/�/??? (?:?L?^?t?�?�?�?l�?��S_�RE�p�d�utLEX$e�[�1-e/VM�PHASE  �!%qCܲxqOFF���_ENB  �<�$VP2��fS�ۯ�@x]#����A@�T����B{�?Gs33������A�m�B�D�Aʼxq� i-���*_>�<r#`�O� �D"?�e�֟������u_�� @�e߀A���<q*���1���9��-�u�_WBj��_�_ ��o=��_�Wa_Vo�_ -o�_�o�o�o�o oco�o;o0Bqoc �oo���o�� %�I[�K�Y�k� ���������3� ُ��1�C�U����� ���ܟ���y�� E�?���~�����џƯ ���Q�����-�s� h���������߯��;� ݿ��+�]���-ϓ� �Ϛ�ɿ��%������� 5�*�Y�K�}�rߡϳπ�ϣ߱�������QTD_FILTE� �j!+ ��& �Ȃ�I�[�m���� ��������C�3��*� <�N�`�r����������	)SHIFTME�NU 1k�-<�<%�?�4��U ,>�bt��� �	��?(u�L	LIVE/�SNAPivs�fliv4N��� ION l@U<��menu��@_$/6/�����ClY����MO�Cm N��zQWAITDINEND  D%��Ai"�&OKsH�/O�UT�/�(S�/�)T�IM�%��	<G �/+=�/N;�/.:�/.:<?�(RELEKAtKf�(TMz;e$��#_ACT�sH'A�(�_DATA n�U(B%8/^O��BR�DIS��>�$�XVRW!o.��$ZABC_GRoP 1pUQ� ,e�2fO��Z�D6@CSCHY q�?I�!���KIPV"r�K%�h�__q_�_�I�MPCF_G 1s�I� P0Rf��_d�Y�Ct�IPpS�� 	�_$o  �<�  ?��  ���;4��aѿB`���DIa4��QaC�����
B׆�>a�>a�C���?����� � \��?�?C��-o?o Qocouo�o�m:�	'o�oNa� ���C��F���������=�?	Y=�Jewx ^x�a�������o�o�o�b0�o�o�D�PY u:_v�_CY�LIND�v�[� �:� ,(  *ȏٍA�ŏ��&�� ?\�n��� ���ǟ������@� !�3�E���i��꟟� ��ï������n��Bs2w�G*A ��_ V���;��7����F���:ז��A���S�PHERE 2x���]�9ϭ�2�o�V� ��ۯ�����W��Ϟ� ��5��Y�@߲Ϗߡ� ������J�������1�`x�U�g�y�@ZZ�6 �e&