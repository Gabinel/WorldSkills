��   b�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����CELLSET_�T   w�$GI_STYS�EL_P �7T  7I�SO:iRibDiTRA�R��I_INI; ����bU9ART�aRSRPNS1TQ234U5678Q�
TROBQACKSNO�� )�7�E�S��a�o�z2� 3 4 5 6� 7 8awn&GINm'D�&��)% ��)4%��)P%��)fl%SN�{(OU���!7� OPTNA �73�73.:B<;}Ta6.:C<;CK;CaI_DECSNAp�3R�3�TRY1���4��4�PTH�CN�8D�D�INCYC@HG�KD~�TASKOK� {D�{D�7:�E�U: �Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T�8�T�@REQ�d��drG�:Mf�GJO?_HFAUL�Xd8�dvgALE� �g�c�g�cvgE� �H�dvgNDBR�H�dg�RGAB�XtbL��c�CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  �0�}qIRTUAALi{q'61�r���p��q�t+ U�P0 �xS�tyle Select 	  ����r�uReq. /�Echo���A�ck���Initiat�p�r�E
�^�m����ʠ�	��
��  ���������������χ�q)��O�ption biGt A<��p�B���C4�Decis��codY��Tr?yout mj�6��Path seg�h�ntin.8�I�g�ycX�:�Tas�k OK?�Ma�nual optK.r�A���B����C� decs�n ��$�Robo�t interl�o7�@�\� iso)lQ�4�C��iM�@���ment<�)��������Ě}�stat�us=�	MH F�ault:����Aler�1�C��p@r7 1�z j�;��y���I�; LE_COMNT ?�y�   Չ�ѿ �����*�<�N�`� rυϖϨϺ������� ��&�9�J�\�n߀� �ߤ߶����������"�����U��Ђ��Ŵ�   ��ENAB  ��:��������������ꮵME�NU\��y��NAM�E ?%��(%$*R�זb��P���t� ��������������+ O:s^p�� ���� $ 6HZ�~��� ����/ /Y/D/ }/h/�/�/�/�/�/�/ �/?
?C?.?@?R?d? v?�?�?�?�?�?�?�? OM