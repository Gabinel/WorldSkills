��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� �~�0COUPLE, �  $�!PP�V1CES C G1��!�PR0�2	 �� $SOFT��T_IDBTO�TAL_EQ� �Q1]@NO`BU SP?I_INDE]uE�XBSCREENu_�4BSIG�0�O%KW@PK_�FI0	$T�HKY�GPANE�hD � DUMM�Y1d�D�!U4� Q �ARG1R��
 � $TIT1d ��� 7T@d7T� 7TP7T55VU65V75V85V95W05W>W�A7URWQ7U�fW1pW1zW1�W1��W 6P!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1�UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t��d�MO� �sE' � [M�s���2�REV�BI�LF��1XI� %�R�  � OD�}`j�$NO`M�+��b�x�/�"u�� ����Q�X�@Dd p =E RD_Eb��?$FSSB�&W`�KBD_SE2uAUG� G�2 "_��B�� V�t:5`ׁ8QC �a_EDu �� � C2�2�`S�p�4%$l �tO$OP�@QB�q�y�_OK���0, P_C� y��dh�U �`/LACI�!�a��x�� FqCOMM� �0$D��ϑ�@�p�X��ORB�IGALwLOW� (KtD2�2�@VAR5�0d!�AB e`BL[@S � ,KJqM�H`9S�pZ@M_O]z�ޗ�CFd �X�0GR@��M�NFLI���;@UIRE�84�"� �SWIT=$/0_NZo`S�"CFd0M�� �#PEED��!�%`���p3`%J3tV�&$E�.�.p`L��ELBOF� �m��m�p/0$��CP�� F�B�����1��r@1J1E-_y_T>!Բ�`���g���G� }�0WARNMxp��d�%`�V`NST�� COR-rF�LTR�TRAT� T�`� $AC�CqM�� R�r$�ORI�.&ӧRT��SFg CHG*V0I�p�T��PA*�I{�T�P�|�� � �#8@a���HDR�B�ą2�BJ; �C��3��4�5�6�7
�8�9>���x@�2� @� TRQB��$%f��ր���֣_U���ѡ�Oc <� ����Ȩ3��2��LLECM�>-�MULTIV4�"�$��A
2q�CHILaD>�
1��z@T_1b�  4� STAY2�b4�=@�)2�4����=�� A|9$��T�A�I`��E��eTO���E��EXT���ᗑ�B��22�0>��@��1b.'��}!9�A�K�  �"K� /%�a��R���?s!>�O�!M��;A�֗�M8�� 	�  =�I�" L�0[�� �R�pA��$JOB�B������TRIGI�# dӀ�����R�-'r��A�ҧ��_�M��b$ tӀF�L6�BNG�A��TBA� ϑ�!��
/1��À�0���R0�P�/p ����%�@|��Bq@W�
2JW�S_RH�CZJZ�T_zJ?�D/5C�@	�ӧ��@����Rd&������ȯ�q�GӨg@NHANC��$LG/��a2qӐ� ـ@��A�p� ���aR��>$x��?#3DB�?#RA�c?#AZt@�(.�����`gFCT����_F�L�`�SM��!I�+ lA�%` �` ���$ /�/����[�a���M�0\��`��أHK���AEs@͐�!�"WꍠN� SbXYZ�W�`�"����6	�������'  �. II��2�(p�STD_C�t�1Q��WUSTڒU�)#�j0U[�%?IO1���� _Up�q�*c \��=�#AORzs 8Bp;�]��`O6  RSY�G�0�q^EUp���H`G�� ��]�DB�PXWORK�+~* $SKP_�p���DB�TR�p , �=�`����Z m�OD3��a _�C"�;b�C� �GPL :c�a�tőS�D�W�3Bb����P�6.� )DB�!��-�B APR��
���DJa3��. p/�u����� �LuYI/�_����0�_^���PC�1�_�S~�EG�]� 2��_�SVPRE.��R3�H $C��7.$L8c/$uSނ�z IkINE�WA_D1%�ROyp��ŀ����q�c7 t@�fP�A���RETUR�N�b�MMR"U���I�CRg`EWM�@�SIGNZ�A� ���e� 0{$P'�1$P� &m�2p�p'tm�+pD�@ �'�bdNa|)r�GO_AW ���@ؑB1I�CYSd�(�CYI�4��B�`1w�qu��t2�z2�vN�}��E}s�DEVIs` 5� P $��RB���I�wPk��IG_BY���"�T7Q��tHNDG�Q6� H4��1�w��$DSBLC��o��v�g@��sPqL��70O�f@]���FB���FEra8�ׂ�t}s��
�8> i�T1?���MCS���fD �ւ
[2H� W��EE����%F����t����9 �T�p��x�NK_N�:�����U��L�wH%A�vZ' ~�2��p�P~r�q7: �='MDLn���9�ጂ ٱh����!e����J��~�+����,�N�D����3��ՒG�!aqSLAd�7;;  ��INP��"�`����}q_ �4<�0�6`C� NU���  D�Lק��S)H!�7=M��q���ܢӢ���g�~��>P +$ٰ �٢��^��^�Y�FI B\��Ă���'A	'AWl�NT�V��]�V~�X�SKI�#T���a�ۺӒT1J�3:3_�P�S�AFN���_SV>�EXCLU��N@��DV@Ll @�Yx����S�HI_V
0^\2PPLYPRo��HIM�T�n�_ML�X��pVRFY_t�Cl�M��IOC�UC_� ����O��q�LS�0M2FT4�Q�����@P҄E$�t��A��CNFK66եu��pm�4ACHD�o�������AFC CPlV�T�QTP?�� �� ?�`�@TA�@�0L@� ��N��]� I@����T��T! S�����te@{RA D8O�� w2���!n��_1�#�HP!�̔�΀K��B�2���MARGI�$����A ��_SkGNE�C;
$ �`�a^aR0��3��@ �B��B��ANNUN�P?���uCN@�`%0����� ����BEFc@I�RD �@Q�F���4OT �`�sFT�HR,Q��CQZ0�M��NI|RE��ȃ���AW���DA=Y=CLOAD�t;T�|�<S5}�EFF_WAXI��F`1Q�O3O��Eq��@_�RTRQE�G�����0RQj�Evp ���F�0f�R�0 �tm�AMP��E<� H 0��`œ^�`Ds�DiU�`���BCAr�' I?�`N Er�IDLE_PWR�I\V!n0V�wV_�[ ꐅ �DIAG��5J� 1$V�`SE�3TQl��e��Pl�^E_l��j�VE� �0SWH�q(� �b2�Gn�OHx3PPHk�IRAl�B�@�[��a�bk�� �w3�O � ��v���I�0 �pRQ�DW�MS-�%A�X{6j�LIFE �@�&�MQy�NH!�Q%��F#C����C(B0�mpN$�Y @�agFLAl���OV0�]&HE��l�SUP�PO�@L1y��@_�$��!_X83�$gq
�'Z�*W�*B1�'T��#`�k2XZáj�Y2D8CY`T@�`!N����f� �C��k���ICTA�K{ `�pCACH��@��3����I��bNӰoUFFI� \� �@��;T��<S6CQBwMSW�5L 8	�KEYIMAG�cTMLa��*Ax�&E��|�B��OCVIER�-aM ��BGLx����y�?� 	��ԣП4N�:�ST�!�BP�D,P�D���D��@EMAI�䐔a��m�r�FAUL|RObB�c�� "spUʰMA"`T'`E�?P< $S��S[ � ITw�BU!F�7y��7�tN[�L'SUB1T�Cx�o�8R�tRSAV|U>R�'c2�\�WT���P �T�*`Sn�_1PbU����YOT�bK��P«�M��d���WAX���2��X1P��S_uGH#
M�YN_�.��Q <Q�D��0����M�� T��F�`|�\�DI��EDT_Pɰ:�IR��b�GRQM�&��HJq�a���׀��Fs�� S (�SV qpB��4�_���a��?T� �@����B�SC_R]1IK >B'r��$t��R"A#u��H�aDSP:FrP�lyIM|Sas�qzՄ�a� U>w� <1%sM�@IP��s��0`tCTHb0ЃTr��T`�asHS�cCsBSCʴq0� V�����S��_D��CONV�E�G���b0^v1PF�Hy�dCs�`&a?ASqC���sMERg�>�aFBCMPg��`�ET[� UBFMU� DU%P�D�:12�CDWy�p�P�C�G�[@NO6�:�V � ��� ���P���EC�����w��A���`��WH *�LƠ�Cc�W���� Y�賂��р�q�|񠀖��A��7}�8B}�9}�H ���1��U1��1��1��1ʚU1ך1�1�2���2����2��2��2���2ʚ2ך2�2*�3��3��3����U3��3��3ʚ3ך�3�3�4��QEXT[�X[b�H``@t&``z�k`˷$����FDR�YTPV��RK"	��K"�REM*F��]"O�VM:s/�A8�TR�OV8�DT�PX�MXg�IN8ɉ W��'INDv�["
�ȕ`K ^`G1a�a��@Q%r7Da�RIV���u"]"GEAR:qI%O.K(�[$N�`����,(�F@� \#Z_�MCM<0K! �Fr� UT���Z ,��TQ? b�y@\t�G?t�E �|�q>Q����[ j�Pa� RI�E���UP2_ 3\ �@=STD	p<TT���������a>RwBACUb] T��>R�d)�j%C�E��0��IFI��0��i��{�4�PTT��FL{UI�D^ �?0gHPUR�gQ�"�r��a�4P+ I�$���Sd�?x��J�`CO�P�SVRT|��N�x$SHO* ��CASS��Qw%�pٴBG_%��3�����FO�RC�B��o�DAT�A��_�BFU_�1��bb�2�en�b0��`� |��NAV	`S������$�S�B~u#$VISI��6�2SC	dSE����j�V��O�$&��BK�� ��$P�O��I��F�MR2��a ��	��`#ǀ�&�8�O� (�_r����+IT_^��ۄ)M�����DG�CLF�DGDY&�LD����5Y&�ϤQ$Y�M됇CbN@~{	 T�FS�P�Dc P��W�cK $EX_WnW�1%`]��"X3�5��G+�d ����SWeUO�D�EBUG��-�G�R��;@U�BKUv��O1R� _ PO_ )������M��LOOc>!S�M� E�R�a��u _?E e >@�G�TERM`%f>i'�ORI�ae 9gi&�`SM_�`>RBe hi%V�(ii%�3UP\Bj� -���e��w#� �f��G�*ELT�O�A�bF�FIG��2�a_���@�$�$g�$UFR�b$`�1R0օ� OT_7�F�TA�p q3NST�`PAT�q�0�2OPTHJ�ԀE�@:�c3ART�P'5p�Q�B�aREL�:�aSHFT�r�a�1��8_��R��у�& � $�'@i�
�����s@bSHI�0�Uzy� �QAYLO�p �Oaq�����1����pERV��XA��H ��m7�`�2%�P�E3��P�RC���ASY1M�a��aWJ07�����E�ӷ1�I��ׁU�T�`Oa�5�F�5P��su@J�7FOR�`MF  �O!k]���5&�0L0���HOL ;l �s2T����OC1!E�$OP��qn���#$�����$��P�R^��aOU��3e��R�5e�X�1 ��e$PWR��IMe�BR_�S�4�� �3�aUD���`�Q�d]m��$H�e!�`�ADDR˶HR!GP�2�a�a�a ��R��.[�n H��S����%��e3��e���e��S�E��L�HS�MNu�o���P��q��0OL�s߰`xڵ�I ACRO��<&1��ND_C�s�x�AfdK�ROUP�B�R_�В� �Q1|� =�s���y%��y-��x@���y���y>�=A��<Ҁ�AVED�w-���u�`(qp $���P_D�� ��'r�PRM_��H�TTP_�H[�q; (ÀOBJ��b6 �$˶LE~3�P|��\�r � ����ྰ_��TE#ԂS��PIC��KRLPiHITCOU�!��L���PԂ������P�R��PSSB�{�JQ�UERY_FLA�vs�@_WEBSOC���HW�#1���s�`<PINCP	U(���O���g������d��t��O���IOLN�t 8�R��$SL�!$INPUTM_U!$`��PLw�֐SL.���u���2�.��C��B�{IOa�F_AS=v�$L+ਇ+�A��bb41�����Z@HYʷ����#q�e�UOP:w ` v�ϡ˶�¡�������"`PIC`���� �|	�H�IP_ME��nv�x Xv�IP�`(�R�_N�p�d����Rʳp�ױQrSP0 �z�C��BG(� r��M�Av�y lv�@CTApB��AL T�I�3UfP_ ۵�0PmSڶBU_ ID�  
�L � `�a�����&0z)����ϴ��NN�_ O��IR�CA_CNf� �{ �Ɖ-�CYpEA��������IC�ǫ�tpR�=QD�AY_
��NTVA�����!��5����gSCAj@��CL�D
����
���v�|5ϰVĬ2b�l�N_�PC V�n�
���w�})�T� �S�����
��e���~T� 2| $Ą �v�~��֣�ذL�AB1��_ ��UN�IX��ӑ ITY裪��ea�R� ��<�)���R_URLn���$A;qEN ����s`vsTeqT_�U���J��X�M�$���E�ᒐR�祪�� A�,���J�H���FLy��= 
|���
�UJR|U� ���F�6G���K7��D>�$J7,�s��J8*�7���$3�E�7��&�8\�)�oAPHIQ4�zy�DkJ7J8Rޒ�L_KE'� o �K͐LMX�� � <U�XR�i�����WATCH�_VAZqu@AំF'IEL`��cyn���&:� � u1VbwP�CTX�j����LGE���� !��LG_SIZ΄�[8Zm�ZFDeIYp1! gXb ZW �S`� 8�m��� �b ���A�0_i0_CM c3#�*'FQ1�KW d(V(Bbpo pm�p� |Io�1 pb p�W RS��0  M(C�LN�R�۠-�DE6E3��� �c�i���PL#�7DAU"%EAq�͐�T8". GH�R��y��BOO�a��3 C��F�ITV�l$�A0��RE���(SCRX����D&�ǒ�qMARGI4�Sp�,@����T�"�y�S���x�W�$y�$��JG=M7MNCHt�y�FN��6K@7r�>9�UFL87@L8FWDvL8HL�9STPL:�VL8"�L8s L8RS"�9HOPh;��C9D�3 R��}P�'IUh�`4@�'�5$ ��S2G09�pPOWG�:�%�3,�64��N9EX��TUI>5I� �ӌ���� �C3�C<0'�,�o�:��&�@�!NaqvcAcNAy��Q�AI]�8gt7Ӝ�DCS���c�RS�cRROXXOdWS��ÂRoXS{X�(IGNp 
Ђ=10 ��[T�DEV�7LL��HY"*�C �	 8�Tr$f/蛒����3-A�a�	 W�萴��Oqs�S1Je2�Je3Ja��BSPC �# �ƋG`-T��% ��Q�T�r@�&E�f+ST�R9 YBr�a� �$E�fC �k�g��f	v9�CB� L����� ��u� xs뀔�g�q�jt��!^�#_ ���ʐ�v�#Ӡ �s �MC��� ���CL�DP᠜�TRQLaI ���y�tFL���rQ��s5�D���w~��LD�u�t�uORG���1�RESERV��M���M�Œ�t~��� � 	�u�5�t�uSV��p���	1�����RCLMC��M�_�ωА��_C�MDBGh��I����$DEBUGMAS������JU�$T8P��EF�d��pFRQҤߏ � K	HR/S_RU4�bq��yA��$EFREQ6�u!$0YOVEAR�k��f�PU17EFI�%Gq��� �
Y�z�� \8����E�$U�`��g?��
�PSI`
��	��CA ��ʲ��σUY�%�?( �	��MISC�味 d��aRQ��	f��TB� � ���A��AX��𑧪�EXCESg�9d�)M�H�9�u����}qd�SC�` � H�х�_�����P������pKE���+�� &�B_, FL�ICBtB� QUI[RE CMOt�O���얩qLdpMD� ��p{!��5b���?$L�MND!��BI����L �D;>
$INAUT�!
$GRSM�ȧPN�b��C���PST�LH� 4U�LO�C�fRI"��eEX���ANG.R.���O[DA]��q��� �RMF0����i�cr�@mu���$�SU�Piu��FX��IG}G! � ��� cs�F�cs
Fct��ޒ �b5��`E��`T�5�tC��g�TI��7 ;�r�M���� t�MD���)��XP���ԁ��H��.���DIAa��Ӻ�W�!��0aTf���D@#)֡O��ܥ���� �CUBp V	���.���O�!9_��� �{`�c������� |�P�|��0� ��P{�KE8B��e-$B��o�=pND2ւ����2�_TXltXTRAhXS������LO: b����}�L����C�.�&�[�RR}2h��� -��!A�� d$C'ALI���GFQj��2F`RINbn�<;$Rx�SW0ۄ����ABC��D_Jp��{�q��_J3��
��1SP, �q�	P����3��H�9pq��#J�3n���O��QIM耯�CSKAP�zb7?SbJ+���Qb�y�����_AZ��/�ELx�Q.ցOCMP����� RTE�� �c1�0 ���1�t�@ ZSMG�0�Э�JG�pSCL<ʠ��SPH_�P�гf��q�u�RT�ER��n�Pk�_EP�q�`A� �c���DI�Q23U�dDF  ���L�W�VEL�qIN8xr�@�_BLXP.��Y/�J��'$F"pIN���]�C�H9%�".�8!6p_T� �F%a"���^$b��k)�~pDHʠt��\�9`$Vw��_�A$=��~�6&A$��S�h���H �$BE�L� m��_ACC�E� 	8�0I�RC_�q�@�NyT��c$PSʠ
�rL���M4�s9  .7��GP/6��9�7$3"�73S2T�͡_Ga�"�0�1��8�1_MG�}�DD�1�~�FW��p��3�5$32�8D}EKPPABN[7ROgEE�2KaBO��p�Ka��1��$USE_v�SP.��CTRTY4@� Z�� <qYNg�A�@�FR �ѢAM:�N�=R��0O�v1�DINC (��B�4���GY��ENC�L��.�K1X2��H0IN�bIS2�8U��ONT�%N�T23_�~�fSL!O�~�|P��Iذ~� �V�~�$��hpU#�yCQ MVMOSI�1�<�[�1����PER�CH  �S���  �W���SlщR��l�� ��E�0�0PAS2EeL�DP7�ONUЉZ��f�VTRK�RqAY"�?c��aS2�e�c������BP�MOM �B���C�H�}�Cj�a�c�3gBT�DUX ��2S_BCKLSH_CS2Fu:��V����C-�esRoz�A�CLALMJT@��`� ��uCHKe ����GLRTYpн�8T���5���_�ùT_UM3��vC3��1Z���7LMT��_LG��%���0�E*�K�=�)� @5F�@8 9�Nb��)hPC�Q)hHТ��5��uCMC���0�7C�N_��N���;S	F�!iV�B��.W�p��S2/�ĈCAT�~SH�Å��4 V�q/q�/V�T1��0PAL�t�B_P�u�c_f �Z�f�Pe�cݔ�uJaG���ѓ�OGއ>�TORQU~@ �S�i @e��R� @B�_Wu�d�!a��#�`��#`�Ih�Iv�I�#F��S�:��I�0�VC00��֢1�ܮ�0��JRK�ܬ!��<�DBXMtt�<�M�_DL�!_bGRVg�`��#`��#A�H_%�?��0���COS��� ��LN #���ߥŴ� ��=�� ����꼰�<�Z���VA�MYǱ:ȧ��᯻�[�THET0�UN�K23�#���#ȰC�B��CB�#Cz�AS�ѯ����#�����SB�#��GTSkZAC����&<���$DU�phg�6�j��E�%Q%a_���x�NEhs1K �t�� y�A}Ŧ�p�׍�����LPH����^U��Sߥ����Ӏ�����!��(Ʀ�V���V�غ ��V��V���V
�V�V&�V
4�VB�H�������ݨd�����H
�H�H�&�H4�HB�O��OR��Os���O��O��UO
�O�O&�O4�O(�F�Ҫ�	����SPBALANgCE_J�6LE��H_}�SP>!۶^��^��PFULC�b�q���K*1��UTO_�p�uTg1T2�	
22N�q 2VP�M�a� i�Z23	qTu`O�1Q��INSEG2�QR�EV�PGQDIF̞ep)1�U�1���`OBK�qj�w2�,�VP�qI�LCHW3AR4B�BAB��u?$MECH��J�X�A��vAX�aPo�p��׫"� � 
��?�10UROB�PCaRS2#%Ղ�@�C1�_ɒT � x� $WEIGH��@�`$��\#��I̾A�PIFvA�0LA�G�B��S�B:�BBIL�%OD�`�Ps"ST0s"P:�pt �� N�C!L �P 
�P2�Aɑ  2���Tx&DEBU�#L�|0�"5�MMY9�C59N��$4�`$D|1 a$0ېl�w > DO_:0AK!� <_ �&� H�q�A��B�"� NJSR�8_�P�@��"O�p �� %�T7P?Q�TL4F0�TICK�#�T1"N0%�3=p�0N�P� u3�PR\p�A��5�|�5U0PROMP�C�E�� $IR�"��A�p8BX`wBMA�IF��A�BQE_� �OCX�a�@RU�C�OD�#FU�@�&I�D_�P�E82B> G�_SUFF�� ��#�AXA�2DO`�7/�5� �6GR�# ��DC�D��E��EP-��DU4� �_ H�_FI�!9GSO�RD�! R 23�6s�HR�AN0$Z�DT�E�`�!X5��4 *WL_NA��1�0�R�5DEF_I�X�RF�T�5�"�6��$�6�S�5�UFIS�m�#�m1|��40c�3��T6�44􁆂�"DP� ?rfd�#D�O@ >l2LOCKE���C��?OG2a�B�@UM �E�R�D�S�D�U�D>b �B�c�E�S�Dd�B�& 2v2a�C�ʑ�E�R�E@�S�C9wwu�H�0P}  d�0,a��F0W�h�u��c=!TE�qY4�� �!LOM�B_�r�w0s"VI]S��ITYs"Aۑ}O�#A_FRI���~SI,a�n�R��07��07�3�#s"WB�W�Q��%�_���AEAS{#�B��P|�x`WB8�45�55��6|#ORMULA�_I���G�W�� h 
>75C?OEFF_O�1&H)��1��Go�{#S� �52CA� :?L3�!G�Rm� � � �$�`�v2X�0TM�g���e�2�c��3�ERIT�d�T� ��  �LL�Dp`SΛ�_SVkd��$��v� �.���� � ���SETU,cMEAG@�@Πt �!HR>L � � (�  0��l��l��aDw��R�0�a�a}d�]�d��B��Ay`�Gax`��[Ѐk@R�EC[Qq�R0MS�K_A y�� P~_!1_USER������*���VE�L����-�!��I�zPB�MT�1CF}G���  �0z]O�NOREJ �0l���[�� �4 e���"�XYZ<SB� 3:!��o_ERRK!� U ѐ�1�@c�Ȱ�!��>�B0BUFIN�DX��R0� MORny�� H_ CUȱ �1��dAyQ?�I>QO$ +�aМ���� \�G{�� ?� $SI�h��@2	�VOv�q�- �OBJE| w�ADcJUF2yĈ�AY��4���D��OUKP�����AMR=�T���-���X2DIR�����Xf�1  DY�Nt�0�-�T� ��R���0� ���OPW�OR�� �,>B0SYSBU�����SOPo���z�U�y�XP�`K���PA`�q������OP�@U���}�"1��/IMAG۱_ ��f�"IM.���IN�������RGOVRD"ё�	���P����  �>gplcC��L�`B�Ű?l�PMC_E(�P�1N��Mr�1b212R�"�SL| ���� �R OVSuL=S�rDEX\aD`��2�:�_"� ��P#���P������2�C �P>���^#�_ZERl���:���� @��:��MO�@RIy��
[�`g@e���s�P�PL����  $FR+EEY�EU�~�Z*��L����T�� �ATUSk�,1C_T�����B�������p�Vc1��P��� !Dc1�к���LQ��`��MQ��ۡL�XE�� x�5IP�W�` ���UP��H`&aPX�;@��43�����PGY��g�$SUB���q���JMPWAIT~ ���LOW���1w�� CVF_A�0���R�Z��CC �R�$��28IGNR_{PL��DBTB� P*a�BW@.t��U�0-IG��!@I��TNLN,�R�Bѡb�N!@��PE�ED~ ��HADO!W� ��t���E�������PSPD��� L_ A�нP��Æ	#UNq � �R�P (�LYwPa�����PH_PK���~b�RETRIE���x���2�R!D@FI���� ���V �$ �2�d�DBGL�V<LOGSIZ,z�baKTU���$�D��_TXV�E�M�Cڡ)�� �-R��#�r��CHECK�z����L���ϰ�q)�L��NPAB�`TJ"����)1P����
�AR�"�BC �=Sa��O�@����ATTS�u䡳&� w�^a�3-#UX^�4�sPL�@Z�� $d�~�qSWITCH�Zh�W��AS��f��3LLB���_ $BA�Dvc��BAMi��6I��(@J5��N�UB6|[F
A_KNOWK34qB"�U��AD+Hc�� D��IPAYL#OAq�9p�C_���GTrѼGZ�CLqAj���PLCL_6� !4��BOA?�T7�VFYCӐ�Jp��D�I�HRՐ�G粒TB��6�J(�zQ_�J�A �B�AND�����T�BQ�q��P�L@AL_ �@�0 =�TAe��pC��uD�CE���J3�P��V� T�PDC�K^�)b��COM�_�ALPH�ScBE0<�߁�_�\�X�x>\� � ���OWD_1�J2�DDM�AR<�h�e�f�cQѯTIA4�i5�i6��MOM(��c�c�ch�c�cV�B� AD�cpv�cv�cPUBP�R�d<u�c<u�b}"�1����� L$PI$��pc��G�y�T�I�yI�{I�{I�s��`�A���v��v��J�b��a��HIG�3���0��� 5�0�f�?�5N�5�SAMPD Ƣ��0����;@�S  ��с6���1���� � ��`���`1�K�P��`�腽P�H��IN 1��P��8�T�/��:��z�Q�z���GAMM�&�S��$GE�T�����D^d>�
�$�PIBR��I.��$HI��_���$1��E=��A�9�*�LW�W�N�9�{��*�Zb���QCdC�HK0�j�ݠnI_��M�JļRoh�Q ���sJ�-v��S ��$�X 1��N�I�RCH_D$RN���^�LE��i�p�Zh8�}ţMSWFL/�M�PSCR�75�Ҽ ��3�"Ķ�6���`��ع�紙��0SV��P'�������GRO�g�S_�SA=AH�=ńNO^`Ci�_d=��no �O�O�x�ʚ��p�B�u,�ȐcDO�A��! �ں�*�t�:�Z1f��;�7����CFMmu�o � �YL�snQ ��� ���"��<s�	�����nQ�8��<3M_Wl���A��\p��(�o�MC ��P���Q���ȇ�hpM.�pr� !��!��$�WM��ANGL�!�AM�6d K�=dK�DdK��TT7�ANk@��3�#�PXC 	OEc�QZ��hp	nt�� ���OM� ��ϑϣϵ����`� �c�Z0es^a_�2� |a�J��i���c�� �cJ��j�����jA畏  � z����  �@{�P�1�P�MON_QU�� �� 860QCO�U��QTHxH�O��B HYS�0ESPBB UE- 3�f0]O�4�  c P��^�RUN_TOʹ�I�O��� �P�@��IND9E�#_PGRA���0���2��NE_NO���ITf��o INFO��a"��ژ��H�OI� =(*�SLEQ!�*0�*�Q OS��l4�� 460ENA�By� PTION��3��r��^GC]F�!� @60J�,�Q���R�d!���erPEDITN�� �� ��KAQj"� �E(�NU'�(AUTY�%CO�PYAQ�2,�qe�M��N< @+��PRU�Tm� C"N�OU��2$G��$R�GADJ��u2X_��IX����&���&W�(P�(~��&9�� z
�N�P_CYCy�e1RGNSc֜{�s�LGO£�NYQ_FREQSrAW@��X1�4�L�@��2P0�!�c@�"�CR1E��MàIF�q��NA��%�4_G>f�STATU~�f���MAIL��|CI<q�=LAST�1a�*4ELEMg� ���QrFEASI t;�ւΰ��B"�F�AF����I� ��O2`�E u�vBAB��PE� =�VA�FzQ��I��TqU[��R���S�FRMS_TRpC�Qc��C��Z�
���1�D I�,2ns�؆�	MB 2� `���N�3V�R2W R*���шR^W�wj�'DOU�^�N�,2�PR`�h�1GR�ID��BARSF!�TYuZ�Op��� |_�4!�� �R�TO��d� � ����PORp�c~vbSRV�0Y)"dfDI[�T�`@;aNd�pXg
�Xg4ViT��Xg6Vi7Vi8:a�v�Fʒg�z $VALU�C0�3D1A�C�ad�� !pf���S�1-Ȇ#AN/��c�0R�]1>1ATOTAL����=sPWE3I�QStR�EGENQzfr��X��H�]5	v( TR�CS�Qq_S3��wfp��V�!��r��BE��3�PG0B�( sV_H�PDA(��p�GS_Ya���i6S��{AR(�2� �"IG_SE�3�pb��5_� �tC_�V$gCMPl��DEp�)G���IšZ~�X��
��Fm�HANC�.� p Qr8�2���INT9`cq��F���MASK\�3�@OVRMP  �PD�1-��W�QaЂ�T�l�_RF�{�V�OPSLGP�g��9�j5��,�;pDpS8���4��U��.��}�TE���`����`k���J^�Y�y3IL_Mx4�s��p��TQ( ���@����5V.�C<�P_ �R��F�M]�V1\�V1�j�2y�2j�3y�3
j�4y�4j���p۲`������ܲIN�VIB8�6�#��*�U2&�22�3&�32��4&�42��6���S�J�  �T $�MC_FK `�B �L>�J�х1pMj�1Iу��zS ��1������KEEP_H/NADD��!鴓@�C��0	��Q����
�O!�v ���p�
�և
�REM!�@	�Cq�RF�]�b�U�4�e	�HPWD  ;�SBM���P?COLLAB*�ph��/q�2IT/0���Q"NO1�FCAqLp⎵��� , ��FLv�A$SY�N���M��Ck��~RpUP_DLY�=�zDELA9�DqZ�2Y AD(����QSKIPO�� i�`� O��NT����c�P_� ��׾  ��cp���q�ٞ��o` ��|`�ډ`�ږ`�ڣ`�ڰ`��9�!�J2�R0  �lX�@T R3H��1AH� �H�8��PRDCq��W� � R�R, 5��R�1��E��5T�RGE�_C��RF#LG"���W�5T�SPC�1UM_|H��2TH2N}Q��;� 1� ��;��Q02 �� D� ˈ��@2'_PC3W�S���1�Y0L10_Cw2���,��� � $\� U@��V7�� ���0��VU\������� rd��C Q +��7��DZ �Gs�RUVL1[�1�h���10]�_D�S�������PK 11�� lڰ����q��AT?��$�Q[7 �� ��K 5T����HOME� *�c2h�n��X��� _3h����!3E )��c4h�hz0���� y�b5h���	//-/(?/&0`6h�b/t/��/�/�/�/�7h��/�/??'?9?�'8h�\?n?�?�?�?�?�WS����  ��Aa{p�����+�_�Ed� T0=�nD4vnCIO䑎I�I@`�O��_OP��E�C.r��WPOW=E	�� X@��f��$$C�d�S����j@�5�3�3� �@�sSI��GP�0�QIRTU�AL�O
QAAVM_WRK 2 7U� ?0  �5Qn_rzXk_�] �\A	�P�]�_3�8P��_�_�Ve�\#m/o�Q`5ojo|o�dHPBS��� 1Y� <Xo�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯz�bC$�AXLM�@t��R��c  d��IN����PRE�
�E�J�-�_U�P��[�7QHPIO�CNV_�� �	�Pr�US>��g�c{IO)�V 1U[P $E`��Qս9lҿ8P?������� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o��o�m�LARMRECOV a���-���LMDG ���ɰ�LM?_IF ��� ை����zv����%�6�, 
 6�_��r漅�������̍$w���׏���8�J�\�n����NGTOL  a�� 	 A   ���ț�PPINFoO ={ <v�����1��   I�3�a�"rP���t��� �����ί���>�o����j�|������� Ŀֿ�����0�B��PzPPLICAT�ION ?����+��Handling�Tool �� �
V9.30P/�04ǐM�
88g340�å�F0����202�ťʚϬ�7DF3��M̎��NoneM�F{RAM� 6���Z�_ACTIVE��b  sï�  ~p�UTOMODz��A���m�CHGAoPONL�� ���OUPLED 1ey� �������g�CUREQ �1	e{  T�
��	p��w����#r���e�HN���{�HTTHKY��
$r��\[�m���� O�	�'�-�?�Q�c�u� ������������ #);M_q�� ����% 7I[m��� /���/!/3/E/ W/i/{/�/�/�/?�/ �/�/??/?A?S?e? w?�?�?�?O�?�?�? OO+O=OOOaOsO�O �O�O_�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_oo#o5o GoYoko}o�o�o�o�o �o�o1CU gy������ �	��-�?�Q�c���1�TO��|�p�DO_CLEAN��|n��NM  �� �B�T�f�x����%�DSPDRY�R��m�HI���@ /�����,�>�P�b��t���������ίj�MAXa�ۄ��������Xۄ������p�PL�UGG��܇�ӌ�P�RC��B� ���ׯF�OK���ȔSEGF��K������ �.�����,�>�v���LAPӟ澨�� �϶����������"��4�F�X�j߯�TOT�AL�7���USE+NUӰ�� �������1�RGDISPWMMC����C��&��@@Ȓ��Oѐ������_STRI�NG 1
��
��M��Sl��
A�_ITEM1K�  nl�g�y�� �����������	�� -�?�Q�c�u����������I/O S�IGNALE��Tryout M�odeL�Inp���Simulat{edP�OutOVERRА� = 100O�In cycl�P�Prog A�borP���S�tatusN�	H�eartbeat�J�MH Fauyl��Aler�	 ������*8<N` ׃G� ׁY�c����� ////A/S/e/w/�/��/�/�/�/�/�/wWOR��G�-1�?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO8�O�O�NPOE� �@E;�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo�BDEV�Nu`�Obo�o �o�o�o�o�o, >Pbt��������PALT ��E?�A�S�e�w� ��������я���� �+�=�O�a�s����GRI�G뽑1��� ���	��-�?�Q�c� u���������ϯ�� ��)�����R�a� ՟;���������ѿ� ����+�=�O�a�s���ϗϩϻ���O�PREG��y���-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_��q����$ARG_�-0D ?	������� � 	$��	+[��]����������SBN_CONGFIG���� ��CII_S?AVE  ��)����TCELLSETUP ���%  OME_I�O����%MOV�_Hn�����REP�d�����UTOBA�CKY���#��FRA:\�� �����)�'`l ���&� 7"�� 24/0�6{  09:35:24�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� ,,		�����O�G�O __#_%_7_q_[_�_ _�_�_�_�_�_�_%o����D�@TSK � �M&,O��UP3DT�@EGd�`�F�XWZD_ENB8ED��fSTADE��ܖe��XIS�UNOT 2��&�(��� 	 o���G{%��=E��Y�a��pp�U2p�Cp�3p�.p��)p�9Ug~)q{��8� ��=� J6��?o� PDC��k>�G����aME�Tc�2LfE� P� qB+X�BU���B(GB����B�ӺC����}?yPw?���s?Z�@U���?]�@A���}SCRDC�FG 1��. ��z������ԏ�����Q =���H�Z�l�~����� 	�Ɵ-����� �2�`D���域���GR�`��`�O���0NA����	��_ED�C@1n�� 
 ��%-�0EDT�-q����%�p�à�u���������������  ��B��2����*�R�b B���*�q���ϧ���3bϮ�@Ͻϯd?���@��=�O���sϏ�4.� ��{�����W���	����?ߏ�5��j�G�� ��#������}�6��6��Z�����Z� ���I��7��� ��&��λ�&m�������8^ҿ���� 	͇�9K�o��!9*�w��	�S���;��CR ����B/T//�/���w//��РNO_�DEL����GE_�UNUSE���I�GALLOW 1���   (�*SYSTEM�*is	$SER�V_GR�;B0�@REGK5$m3i|B0�NUMp:�3�=P�MU� iuLA�Y�pi|PM�PALD@�5CYC10�.�>�0�>CULSU�?�=�2�A�M3LOWDBOX�ORIt5CUR_�D@�=PMCNV6�6D@10�>�@T4DLI�`=O_9�	*PROGRA�J4PG_MI�>�OPAL�E_U�PB7_B>$F�LUI_RESU`�7p_z?�_�TMRY>h0�,�/�b�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv����������"LAL_OUT 1;�l���WD_ABO�R�0?d�ITR_�RTN  �����g�NONSTO�Ǡ�� 8CE_�RIA_I0���ۀ��ŀFCFG ��۔��o_LIMY22ګ� �  � 	i�J��<e�g��5�� 9���������
���u��P}AQPGP 1�����Q�c�u�b4�CK0����C1���9��@���PC��CUV��]��d��l��as��P���C[٤Um��v�������_�� C����-�m��?�ÂHE� �ONFI�Pq�G�G�_P�@1� �%�������ǿٿ�����G�KPAU�SaA1�ۃ  �2�W��Eσ�iϓ� �ϟ����������#߀I�/�m��eߣ��M~��NFO 1"�;�� �7�������B�J-���]��q9C�����'��f� � �DX��C��Z³��C�+�4�4F�ŀO��c�COLLECT�_�"�[�����E�N�@��y���k�ND-E��"�3�"�1234567890��\1�� �$�֕H&��)M�r� \,L�^���]+������ ������C 2� Vhz���� ��
c.@R��v�������΢� ����IOG !���q���`u/�/�/�/C'TR�K2"'-(׀^)
��.R�#R-�*W� 9�_MOR�$� �;�l5��l9�?r?�?@�?�?�;E2��%S=%,W�?@�@��C׀�K)DցC�R�&�u�XOWAWBC4  �A�q��׀x׀}A"@Cz  B�@�CG�B8��AC [ @yB�׀ց�:d�43 <#�
�E���I�O�C*=AI��'GM?�C��(S=���Qd=AT_�DEFPROG ��;%�/m_APINUSE�V�ۅ�T�KEY_TBL � s�ہ���	
��� !"#�$%&'()*+�,-./�:;<=>?@ABCDP�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������Ga�������������������������������������������������������������$��PL�CK�\���P�PST�An��T_AUTO�_DO��NFsI�ND���n��R_T1wT2N�����5ŀTRLCPLE�TE���z_SCREEN ��kcscÂU���MMENU 1)O� <�[_#� q��,�a���>�d��� t���ӏ����	���� �Q�(�:���^�p��� ����̟�ܟ�;�� $�q�H�Z��������� �Ưد%����4�m� D�V���z���ٿ��¿ �!���
�W�.�@ύ� d�vϜ��ϬϾ���� ��A��*�P߉�`�r� �ߖߨ��������=� �&�s�J�\����������'�,�p_?MANUAL�Eq�DB
12�v�iDB�G_ERRLIP9*�{h! 0��������g�NUML�IM�s:QOE�@D�BPXWORK 1+�{��>Pb�t��-DBTB_��q ,��kC3!�VD!DB_AW�AYo�h!GCP� OB=��A�_A!L���o�k�Y�p�utO@`�_�� 1-�+@
-k-6[�6�_M+pIS�`��@"@�ONTIM6�w�OD��&�
�U;MOTNE�ND�_:RECO�RD 13�{ y��[CG�O�f! T/[K��/�/�/�/_( �/�/f/?�/??Q?c? �/?�??�?,?�?�? OO�?;O�?_O�?�O �O�O�O(O�OLO_pO %_7_I_[_�O_�O�_ _�_�_�_�_l_!o�_ ,o�_io{o�o�oo�o 2o�oVo/A�o eP^�
��� R���=��a�s� �������*�ߏN�� �'���ԏ]�̏���� ����ɟ۟v���n�#����G�Y�k�}���TOLERENC�sB�0� L��g��CSS_CNST_CY 24	�t�	��.������ 0�>�P�b�x������� ��ο����(�:��äDEVICE ;25ӫ ��� �ϱ������������/�AߟģHNDG�D 6ӫ� Cz�T�.!ơLS 27t�S������������/�U�ŢPARAM 8Gb�A���Ք�RBT 2:.8�<����CkA� �~��  � A�p��.SB���~A�B�  ����������.`��  ����A�A�C����c�u����C�A�D��k�epz�A�A��HA�c��A�	�?(u�L^p���A�B�t/�D��C���_ 	 A=���ABffA#�33AҊ��ͳA�A�Cf��aĒ�A�J��7B]���B��B�ffBᴠ�33�C$.@R� ( ����A���� 
/��//)/;/�/ _/q/�/�/�/�/�/�/ �/<??%?r?I?[?m? ?�?�?�?�?�?&O8O �PObOMO�OqO�O�O �O�O�O_�OOL_ #_5_�_Y_k_�_�_�_ �_ o�_�_6ooolo CoUogo�o�o�o�o�o �o �o	h�O� w�����
�� .�	__I'�1_�q� �������ˏݏ�� �%�r�I�[������ ����ǟٟ&����\� 3�E�W����ȯ��� ׯ�"��F�1�j�E� s�����m�������ѿ �0���f�=�O�a� sυϗ��ϻ������ ��'�9�Kߘ�o߁� ����[����(��L� 7�p��m����� ������$�����l� C�U���y��������� �� ��	V-?� cu����
�� @+dO�s� �������*// /`/7/I/[/m//�/ �/�/�/?�/�/?!? 3?E?�?i?{?�?�?�? �?�?�?�?FO�jOUO gO�O�O�O�O�O�O_ _�'O9OO=_O_�_ s_�_�_�_�_�_�_�_ oPo'o9o�o]ooo�o �o�o�o�o�o: #5��O������ ��$��H�Fz��$DCSS_SL�AVE ;����w��~`�_4D  w����AR_MENU <w� >�؏� ��� �2�^rǏ\��n�\���SHOW �2=w� �  fr[q����Ə������,�>�D�b�t���  ����ҟϯ���� )�P�M�_�q������� ��˿ݿ���:�7� I�[ς�|Ϧ��ϵ��� ������$�!�3�E�l� fߐύߟ߱������� ���/�V�P�z�w� ������������ �@�:�d�a�s����� ������\���*�H� N�K]o���� ����28�G Yk}����� �"�1/C/U/g/ y/�/��/�/�/��/ /?-???Q?c?u?�/ �?�?�?�/�??OO )O;OMO_O�?�O�O�O �?�O�?�O__%_7_ I_pOm__�_�O�_�O �_�_�_o!o3oZ_Wo io{o�_�o�_�o�o�o �oDo-Se�o ��o�������.�=�O���CFG7 >�����q���dMC:\���L%04d.C�SV\��pc��������A ՃCH݀z��v�w�#�  ���:�J�8�<S���JP�j�)����p7�-�n�RC_OUT ?z������a�_C_FSI ?��? |�� ���@�;�M�_��� ������Я˯ݯ�� �%�7�`�[�m���� ����ǿ�����8� 3�E�Wπ�{ύϟ��� ���������/�X� S�e�wߠߛ߭߿��� �����0�+�=�O�x� s����������� ��'�P�K�]�o��� ��������������( #5Gpk}�� ��� �H CUg����� ��� //-/?/h/ c/u/�/�/�/�/�/�/ �/??@?;?M?_?�? �?�?�?�?�?�?�?O O%O7O`O[OmOO�O �O�O�O�O�O�O_8_ 3_E_W_�_{_�_�_�_ �_�_�_ooo/oXo Soeowo�o�o�o�o�o �o�o0+=Ox s������� ��'�P�K�]�o��� ��������ۏ���(� #�5�G�p�k�}����� ��şן �����H� C�U�g���������د ӯ��� ��-�?�h� c�u���������Ͽ�� ���@�;�M�_ψ� �ϕϧ���������� �%�7�`�[�m�ߨ� �ߵ����������8� 3�E�W��{����� ���������/�X� S�e�w����������� ����0+=Ox s������ 'PK]o� �������(/ #/5/G/p/k/}/�/�/ �/�/�/ ?�/??H?�C?U3�$DCS_�C_FSO ?�����1? P [?U? �?�?�?�?�?O
OO .OWOROdOvO�O�O�O �O�O�O�O_/_*_<_ N_w_r_�_�_�_�_�_ �_ooo&oOoJo\o no�o�o�o�o�o�o�o �o'"4Foj| �������� �G�B�T�f������� ��׏ҏ�����,� >�g�b�t��������� Ο�����?�:�L� ^���������ϯʯܯ�g?C_RPI~> �?�;�d�_�
�}?.�`p����ݿj>SL�@���9�b�]�oρ� �ϥϷ���������� :�5�G�Y߂�}ߏߡ� �����������1� Z�U�g�y������ ������	�2�-�?�Q� z�u������������� 
)RM_q ������� *%7Irm� ����/�ϛ� ,�/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO sO�O�O�O�O�O�O_ __'_P_K_]_o_�_ �_�_�_�_�_�_�_(o #o5oGopoko}o�o�o �o�o�o �oH CUg��������� ����NOCODE @������PR�E_CHK B쟻3�A 3��< �7�����<���� 	 <��� ��?#ۏ%�7��[�m� G�Y�������ٟ�ş �!����W�i�C��� ��y�ïկˏ���� ��A�S�-�_���c�u� ��ѿ�������=� �)�sυ�_ϩϻϕ� �������'�9���E� o�I�[ߥ߷ߑ����� ����#����Y�k�E� ���{�������� ���C�U��=����� w���������	���� ?Q+u�a�� ����); _qg�Y��S� ���%/�/[/m/ G/�/�/}/�/�/�/�/ ?!?�/E?W?1?c?�? ���?�?o?�?O�? �?AOSO-OwO�OcO�O �O�O�O�O_�O+_=_ _I_s_M___�_�_�_ �_�_�?�_'o9oo]o ooIo�o�oo�o�o�o �o#�oGY3E ��{����� o�C�U��y���e� ����������	��-� ?��K�u�O�a����� ����͟��)��1� _�q��}�������ݯ �ɯ�%���1�[�5� G�����}�ǿٿ��� ����E�W�1�{ύ� G�u����ϯ������ /�A��-�w߉�c߭� �ߙ���������+�=� �a�s�M���ϑ� ������'��3�]� 7�I������������ ������GY3} �i������� �C/y�e �������-/ ?//c/u/O/�/�/�/ �/�/�/�/?)?�? _?q?K?�?�?�?�?�? �?�?O%O�?IO[O5O O�OkO}O�O�O�O�O _�O3_E_;?-_{_�_ '_�_�_�_�_�_�_�_ /oAooeowoQo�o�o �o�o�o�o�o+ 7aW_i_��C� ����'��K�]� 7�i���m��ɏۏ�� �����G�!�3�}� ��i���ş����� �1�C��g�y�S�e� ���������ѯ�-� ��c�u�O������� Ͽ�ןɿ�)�ÿM� _�9�kϕ�oρ����� �������I�#�5� ߑ�kߵ��ߡ����� ��3�E���Q�{�U� g������������ /�	��e�w�Q����� ����������+ Oa�I���� ���K] 7��m���� �/�5/G/!/k/}/ se/�/�/_/�/�/�/ ?1???g?y?S?�? �?�?�?�?�?�?O-O OQOcO=OoO�O�/�/ �O�O{O�O_�O_M_ __9_�_�_o_�_�_�_ �_oo�_7oIo#oUo oYoko�o�o�o�o�o �O�o3Ei{U �������� /�	�S�e�?�Q����� ��я㏽���� O�a�������q���͟ �������9�K�%� W���[�m���ɯ��� ��ٯ�5�+�=�k�}� ������������տ �1��=�g�A�Sϝ� �ω����Ͽ��������Q�c����$D�CS_SGN �CS����#M��24-JU�L-24 12:�22 E�06���N��09:39������� X�L��������������ДќM��?Þ�j������{�VERSION� ��V4�.2.10�EF�LOGIC 1D�S��  	D���X�k�X��z�M�PROG_E_NB  ��b���Л�ULSE  ����M�_AC�CLIM��������WRSTgJNT����w�EMO���ѷ�L��INIT EZ��O��OPT_S�L ?	S�1�
 	R575��V��74��6��7��)5A��1��2��l����G�h�TO  �t���.H�V?�DE�X��d����FP�ATH A��A�\4���HC�P_CLNTID� ?+�b� �l�����IAG_�GRP 2JS�� ��a[�D�  D��� D  B߫  B�@ff��/B�@[���W�@�q���B�N�C�-�Bz��Bp@�e`��mp3�m7 7890123456�*�[���  Ao��mAj1Ad�A]�
AW|��AP�AJ-�AC/A;�ǞA4H���@�W  A��A�A3!�_A�@@��B4�� ��t����
�uƨApf�fAj�yAeK��A_�AY���AS� MC�AF��A@ �O��+/=/O$O�c K�w(@�X?8��@��y�/�/�/�/��/8�;d�2�5�?@~ff@x1�'@q��@kC��@d�D@]��@Vv�6?H?Z?�l?~?8s�0l���@e@^���@W\)@O���@H�0?<@7K�@.V�?�?�?�?|
O8S@M00�G<@A��@<�1@5��@/l�@(Ĝ@!�0�\NO`OrO�O�O x'g�L_K�;_�_�__ g_�_�_�_�_o�_�_ �_YokoIo�o�o+o�oX�"� 2�17A�@�J>��R
q?��33?Y��r{��J7'Ŭ2q�63p4�F>r�{�LJ@�p�Zr��
=@�@��Q�jq��@G A�h�@��@�T= �c<��]>*��H>V>��3�>���J<���<�p�q�x���� �?� ��C�  <(�U��� 4Vr�33���@
���A@��? R�oD��mR�x���Q� �t����Z�Џ��؏��,��i?�7N�>��(�>�@Z�=�{��J��G�v�G�J�B�E�����a���@ǐ@���@~��@Q�?L *���ŲI�PP���&���'���@�K����Ag�q�PC��  C���C!uy�
���ʯ ?�� ��	��Գ�4���X���v���*����DX��C��$³����B�ÿ f��ҿ���A�,�����r>�Ty��H�>~�>� �
�Iϗ��CT_CONFI/G K3��ԟeg��STBF_TTS��
����"��������{�MAU���M_SW_CF��L�  �OCVI�EW	�MI�U��㯛߭߿������� ���0�B�T�f�x� ������������ �,�>�P�b�t���� ������������( :L^p��� ��� �6H Zl~�������/��RCB�N��!��F/{/j/��/�/�/�/�/��SB�L_FAULT �O9*^�1GPM�SK��7��TDI�AG P��U�����qUD�1: 6789012345q2�q���%P�ϭ?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O �a6�I�'�
�?_��TRECPJ?\:
j4\_�7 _[�?�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�O�O_ _��UMP_OPTIcON��>qTRB�t��9;uPME���.Y_TEMP � È�3B�����p�A�pytUN�I'��ŏq6�YN_?BRK Qt�_�?EDITOR q&q�h�r_2PENT �1R9)  ,�&COLOCA�_bpA_IRVI�S$r5� &P�EGA_BARR�A_ESTEIR�A 3���&M�AIN Q���&SEGU��}���P�p��  &�-BCKEDT-� ���pNO��,�&�PROG_1 �׏�SUMIR�P���DROP�_DEFE�p �E#RT:���S�2b�H��Z�3���� �AN?TENA_C���]T�SEMX� 1��� �.����&PICKUP��M����*�(�	���p��ғ(�F��DA_P�RENSA�����\���7�9��\�1?_PLACE0���&
L�4�3�����J�]�.����pMGDI_STA�u�~��q���pNC_I?NFO 1SI��b�������Կ�쮳��1TI� � �o#��P�0�d�o}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������Hu� � 2�D�R�j�R�x��� ������������,� >�P�b�t��������� ����Z��#5G a�k}����� ��1CUg y�������� 	//-/?/Yc/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?��?O%O7O Q/GOmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�? Ooo/o�_[Oeowo �o�o�o�o�o�o�o +=Oas�� ����_�_��'� 9�So]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�K�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�C�5�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� ������!�;�M�W� i�{���������� ����/�A�S�e�w� �������������� +E�Oas�� �����' 9K]o���� 1����/#/=G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?��?�? 	OO5/?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�?�_�_oo-O#o Io[omoo�o�o�o�o �o�o�o!3EW i{����_�_� ���7oA�S�e�w� ��������я���� �+�=�O�a�s����� ����ߟ���/� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������͟׿ ����'�1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߫�ſ�������� �;�M�_�q���� ����������%�7� I�[�m�������߯� �������)�3EW i{������ �/ASew ���������/ !+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?/� �?�?�?�?/#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�?�_�_�_�_ Oo-o?oQocouo�o �o�o�o�o�o�o );M_q���_ ����	o�%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�����ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߩ������� �����1�C�U�g� y������������ 	��-�?�Q�c�u��� �߫����������� );M_q��� ����%7 I[m����� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? ���?�?�?�?�O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�?�?�_�_ �_�_�?�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y�_�����_� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q��y��� ��˟�۟��%�7� I�[�m��������ǯ ٯ����!�3�E�W��i��� �$ENE�TMODE 1U��� + ���������»��RROR_P�ROG %��%������TABL/E  ���Q��c�uσ��SEV_�NUM ��  �������_�AUTO_ENB�  ̵��ݴ_N�O�� V�������  *����J����������+����(�:���FLTR����HIS�Ð������_ALM 1W.�� ����̍�+;����������0�?�_����  ���²u꒰TC�P_VER !�!��@�$EXTLOG_REQv�s�����SIZ����STK��������TOL  ���Dz~��A ��_BWDU�*�Z��V�ǲ?�DID� X�Z�����[�STEPl�~���>��OP_DO����FACTORY_�TUNv�d��DR_GRP 1Y��`�d 	p�.° ��*u����RHB ��2� ��� �e9 ���bt� o��������J5nY@1���A5�@���?ͨeu
? J�9��� uȸo��_/�(/�(B�  F!A���33R"�33^-@UUTn*@�� /ȷ>u.�>*��<��ǆ-�E�� F@ ξ"�5W�%�-J���NJk�I'�PKHu��IP��sF!���-?�  ?�/9��<9�8�96C'6<�,5���-����������,�_s �* &����i$��F�EATURE �Z�V�Ʊ�Handling�Tool �5���English� Diction�ary�74D S�t�0ard�6�5A�nalog I/�O�7�7gle S�hift Outo� Softwar�e Update�%Imatic B�ackup�9SAg�round Ed�it�0�7Came�ra�0F�?Cnr�RndImXC�Lo�mmon cal�ib UI�C�Fn�qA�@Monito�r�Ktr�0Rel�iab@�8DHC�P�IZata A�cquis�CYiagnosOA�1[�ocument �Viewe�BWu�al Check Safety�A~�6hanced�F4�:�UsnPFr�@�7�xt. DIO ��@fiRT�Wend.�PErr�@LQR�]J�Ws�Yr�0�P E���:FCTN Me�nu�Pv S8gTPw In'`facNe�5GigE`nrej@�p Mask Ekxc�Pg�WHT^`�Proxy Sv�oT�figh-Spe�PSki�D�eJP~�PmmunicN@7ons�hurE`'`�_�1abconne�ct 2xncr``stru�2z>p�eeQPJQU�4KA�REL Cmd.� L�`ua�husR�un-Ti�PEnyvkx(`el +R@�sP@S/W�7License�Sn\�P�Book(Sys�tem)�:MAC�ROs,�b/Of'fse@�uH�P8@�_�pMR�@�BP^MechStop�at.p6R�ui�RKj�ax�P�0P@)�od@witch��>�EQy.���OptmЏ�>��`filn\=�g�w�uulti-T��`tC�9PCM funHwF�o3T�R?�^f�Regi�pr�`I�rigPFV����0Num Selb�|���P Adju�`��J�tatu�
�iZ�5RDM �Robot�0scgove�1F�ea7���PFreq An;ly�gRem`��Q�n�7F�R�Serv�o�P���8SNPX� b�rNSN^`C�lifQɮBLibr�3鯢0 q������o�ptE`ssag?��4�� -C��;���/I_mB�MILI�Bk�E�P Fir�m6BU�PEcAcc<k@sKTPTX_C�eln���F��1��V�orqu@imGula�A�A�u���Pa�qU�j@�Ã&ε`ev.B�.@ri�P޿USB poort �@iP�P�agP��R EVN�T�ϗ�nexcept�P��t��ſX�]�VC�Ar�b�bf�V@2PҦ�$����SܠsSCصV�SGEk��a�UI�;Web Pl!��ާ��Խ`��TeQfZDT Appl�d�:�ƺ� ��GridV�pla�y�R�WD4�R
�.��:n�EQ+��r-10�iA/7L*��1G?raphic���5�dv�SDCSJ�c�k�q�5larm �Cause/��e}d�8Ascii�a���LoadnP�U�pl,�Ol�0�AG�u�6N�`���yFyc�@�r�����PV��Jo��m� c�R���c���m�./�����Q�2*u:eRAJ��P�ٌ�4eqinL����8N�RT��9On�0e Hel�HJ�`oI�alletiz?��H�����_�tr�[R?OS Eth�q���T@e�ׅ�!�n�%�2D�tPkg&�Upg~�(2D�V-�3D Tr�i-jQEAưDe�f.qEBa)pde`i��� �bImπqF�f��nsp.q�=�464MB D�RAMZ,#FRO�5/@ell�<�Mshf!r/�'c%3@YpLƖ,ty@s˒xG��m��.[�� ���BU���Q�B�=mai�P߫�]Q����@q6wlu����^`�x�R�?eL� Sup�������0�P�`cr ��@�R���b䚮�pr1ouest�rt~QQ��ߋL!�4O��q�$�K��l Bu�i7�n��APLCdOO�EVl%��CGUN�OCRG�O��DR���O
TLS_��BU�/_��K�qN_d�TA�OxVB�_�W�ܑZ���_TCB�_�V�_�W���WF+o�V�O�W._8�W�ņoTEH�o�f0�O�gt�oTEj�xV!F�_w�_xVGoTw�BTw~oxVH�xVIaA��v�xVLN�yUMz�bo�f_xV	N�xVP���^xV	R&xVS��܇ʏ���W��v���VGF:�L�P2_h��h��V�h��_g�D��h�F0Foh��g�RD�� 7TUT��01:�L�y2V�L�TBGG���v�rain�UI���
%HMI���p#on��m�f�"��F�&KAREL9� �TPj��<6� SWIMEST&ڢF0O�<5�
"a� X�j�������ͿĿֿ ���'��0�]�T�f� �ϊϜ����������� #��,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ ����������$�Q� H�Z���~��������� ���� MDV �z������ 
I@Rv ������// /E/</N/{/r/�/�/ �/�/�/�/???A? 8?J?w?n?�?�?�?�? �?�?O�?O=O4OFO sOjO|O�O�O�O�O�O _�O_9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l���������Ə ����)� �2�_�V� h����������� ��%��.�[�R�d��� ������������!� �*�W�N�`������� �����޿���&� S�J�\ωπϒϤ϶� ��������"�O�F� X߅�|ߎߠ߲����� �����K�B�T�� x����������� ��G�>�P�}�t��� ���������� C:Lyp��� ���	 ?6 Hul~���� �/�/;/2/D/q/ h/z/�/�/�/�/�/? �/
?7?.?@?m?d?v? �?�?�?�?�?�?�?O 3O*O<OiO`OrO�O�O �O�O�O�O�O_/_&_ 8_e_\_n_�_�_�_�_ �_�_�_�_+o"o4oao Xojo|o�o�o�o�o�o �o�o'0]Tf x������� #��,�Y�P�b�t��� ������������ (�U�L�^�p������� ���ܟ���$�Q� H�Z�l�~�������� د��� �M�D�V��h���  �H552}���21n��R78��50���J614��ATU]PͶ545͸6���VCAM��CRIn�UIFͷ28	ƷNRE��52��R�63��SCH��DwOCV]�CSU���869ͷ0ضEI�OC9�4��R69���ESET���J�7��R68��MA{SK��PRXY!�]7��OCO��3�h����̸3�J6˸�53��H2�LCH^��OPLG�0֯MHCR��S{�MkCS�0��55ض�MDSW���OP��MPR�M�@�0n̶PCM �R0���ض��@�51�5u1<�0�PRS�ǻ69�FRD�FwREQ��MCN��{93̶SNBAE�^3�SHLB��M��tM���2̶HTC��TMIL����TP�A��TPTX��EL��Ѐ�8������wJ95,�TUT׻95�UEV��U�EC��UFR�V�CC��O��VIP��CSC,�CSGt8�r�I��WEB�7HTT�R6C�N��CGIG��IP�GS)RC�DG��H77��6ضR�85��R66�Ru7��R:�R530�K680�2�q�J��*H�6<�6,�RJح�j0�4�6o64\��5�NVD��R6��R84Tg�����8�90\���J9&3�91� 7+����,�D0oF�CL9I���CMS�� n�STY��TO䶴q���7�NN�O�RS��J% ��j�O]L(END��L���Sf(FVR��V3�D���PBV,�A�PL��APV�C�CG�CCR|�C�D��CDL@CS�Bt�CSK��CT�CTBL9��U0,(�C��y0L8C��TC� �y0�'TC(7TC���CTE\��07T�Eh��0��TFd8FJ,(GL8GI�8H�8�I��E@�87�CTM�,(M�8M@8N�8P�HHPL8Rd8(TSrd8W�I@VGF�GP2��P2���@�H�{7VPD�HF �V�PSGVPR�&VT���YP��VTB7Vs�IH��VI aH'�VK��VGene�����_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 I[m���� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/?�?+?=?O?a?s?�?�  H55�hT�1�1[U�3R78��<50�9J614έ9ATU�T�454u5�<6�9VCA�Dn�3CRI,KUI8Tv�528-JNRE�:�52JR63�;S{CH�9DOCV�J�CU�4869�;0N�:EIO�TsE4�:�R69JESET��;KJ7KR68ތJMASK�9PR�XYML7�:OCOB\3�<�J)P�<3|Z[J6�<53�JH�\�LCH\ZOPLGz�;0�ZMHCR]Z]SkMCS�<0,[{55�:MDSW}kv�[OP�[MPR�Zt�@�\0�:PCMLJ�R0�k)P�:)`�[5�1K51|0JP�RS[69|ZFR�D<JFREQ�:M�CN�:93�:SN�BA}K�[SHLB��zM�{�@ll2�:H{TC�:TMIL�<��JTPA�JTPT�X�EL�z)`�K8��;�0�JJ95\JT�UT�[95|ZUE�VZUEC\ZUF]R<JVCC��O<jwVIP,�CSC\��CSGlJ�@I�9W�EB�:HTT�:R�6{L��CG{�IG�[�IPGS��RCv,�DG�[H77�<�6�:R85�JR6�6JR7[R|R[53{68|2�ZR�@Jml,|6|6\JQR�\	P|4L�6��64��5�kNVDvZR6+kR84<�h��IP,�8��90��6�KJ9�\91��̫�7[KIP\JD0�F���CLI�lKCMqS�J9��:STY,��TO�:�@�K7�LN]N|ZORS<jJ���MZZ|OLK�END�:L�S��FVR��JV3D,�KKPB�V\�APL�JAP�V�ZCCG�:CC�RjCD�CDL�̚CSB�JCSKv�jCTK�CTB�݈\���\�C�z���C�L�TCLJ�l�TCv��TCZCTE�J���|�TE�J��<�TUF��F\�G��G��
l�Hl�I�z)�l�k�WCTM\�M\�M��UNl�P,�P��R�ܖ;�TS��W��̚V�GF��P2��P2p�z �VPD�FLJVP;�VPR���VT�;� �JVT�B��V�KIH�VXِM�<�VK,�V{�Gene�8�83E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ��������� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ��������1�C�U� g�y������������� ��	-?Qcu ������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ �/�/�/�/?!?3?E?�W?i?{?�7�0�STD�4LANG�4�9�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~��������� �2�D�V�RB=T�6OPTNm�� ������Ǐُ���� !�3�E�W�i�{�����8��ß�5DPN�4� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G��Y�k�}ߏߡ߳�ted �4�8������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u��������� ������);M _q������ �%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ������*�<�N�`�r�99���$F�EAT_ADD �?	�����~��  	�� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu������DEMO �Z��   ���}��'��0� ]�T�f����������� ����#��,�Y�P� b�������������� ���(�U�L�^��� ���������ܯ�� �$�Q�H�Z���~��� �����ؿ��� � M�D�Vσ�zόϦϰ� �������
��I�@� R��v߈ߢ߬����� �����E�<�N�{� r����������� ��A�8�J�w�n��� ������������ =4Fsj|�� ����90 Bofx���� ���/5/,/>/k/ b/t/�/�/�/�/�/�/ �/?1?(?:?g?^?p? �?�?�?�?�?�?�? O -O$O6OcOZOlO�O�O �O�O�O�O�O�O)_ _ 2___V_h_�_�_�_�_ �_�_�_�_%oo.o[o Rodo~o�o�o�o�o�o �o�o!*WN` z������� ��&�S�J�\�v��� �������ڏ��� "�O�F�X�r�|����� ��ߟ֟����K� B�T�n�x�������ۯ ү����G�>�P� j�t�������׿ο� ���C�:�L�f�p� �ϔϦ�������	� � �?�6�H�b�lߙߐ� ������������;� 2�D�^�h������ �������
�7�.�@� Z�d������������� ����3*<V` �������� /&8R\�� �������+/ "/4/N/X/�/|/�/�/ �/�/�/�/�/'??0? J?T?�?x?�?�?�?�? �?�?�?#OO,OFOPO }OtO�O�O�O�O�O�O �O__(_B_L_y_p_ �_�_�_�_�_�_�_o o$o>oHouolo~o�o �o�o�o�o�o  :Dqhz��� ����
��6�@� m�d�v�������ُЏ ����2�<�i�`� r�������՟̟ޟ� ��.�8�e�\�n��� ����ѯȯگ���� *�4�a�X�j������� ͿĿֿ����&�0� ]�T�fϓϊϜ����� �������"�,�Y�P� bߏ߆ߘ��߼����� ����(�U�L�^�� ������������ � �$�Q�H�Z���~��� ������������  MDV�z��� ����I@ Rv����� ��//E/</N/{/ r/�/�/�/�/�/�/�/ 
??A?8?J?w?n?�? �?�?�?�?�?�?OO =O4OFOsOjO|O�O�O �O�O�O�O__9_0_ B_o_f_x_�_�_�_�_ �_�_�_o5o,o>oko boto�o�o�o�o�o�o �o1(:g^p ������� � -�$�6�c�Z�l����� ��ϏƏ؏���)� � 2�_�V�h�������˟ ԟ���%��.�[� R�d�������ǯ��Я ���!��*�W�N�`� ������ÿ��̿�� ��&�S�J�\ωπ� �Ͽ϶��������� "�O�F�X߅�|ߎ߻� �����������K� B�T��x������ �������G�>�P��}�t���������  ������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<N`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz����>�y  �x�q ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^�p������q�p�x���*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p���������������$FEAT_D�EMOIN  V�� �����_INDEX����ILECOM�P [����B��8 S�ETUP2 \�BL�  �N w5_AP2�BCK 1]B	  �)����%����E �	 ���5�Y�f� �B��x/� 1/C/�g/��/�/,/ �/P/�/t/�/?�/?? �/c?u??�?(?�?�? ^?�?�?O)O�?MO�? qO O~O�O6O�OZO�O _�O%_�OI_[_�O_ _�_�_D_�_h_�_�_ 
o3o�_Wo�_{o�oo �o@o�o�ovo�o/ A�oe�o��� N�r���=�� a�s����&���͏\� 񏀏���"�K�ڏo� ������4�ɟX���� ��#���G�Y��}��@��0���ׯQ	� P�� 2� *.V1Rޯ(���*+�Q�`��W�{�e��PC��|����FR6:��"ؾg�����T   � 2����\� ��d��*.F��ϕ�	�ó����o�ߓ�STM�9���ư%�d��ψߓ�HU߻�J���f�x���GIF �A�L�-����ߑ��JPG����Lձ�n������JS�H������6���%
Ja�vaScriptt���CSe���Kֹ��v� %Casc�ading St�yle Shee�ts��j�
ARGNAME.DT'
��O�\;��[�k�|(k DISP*rUOп���� �
TPEIN�S.XML/�:�\CcCust�om Toolb�ar��	PASS�WORD���F�RS:\�� %�Passwor�d Config /c�Q/�J/�/���/ :/�/�/p/?�/)?;? �/_?�/�??$?�?H? �?l?�?O�?7O�?[O mO�?�O O�O�OVO�O zO_�O�OE_�Oi_�O b_�_._�_R_�_�_�_ o�_AoSo�_woo�o *o<o�o`o�o�o�o+ �oO�os��8 ��n��'��� ]�����z���F�ۏ j������5�ďY�k� �������B�T��x� ����C�ҟg����� ��,���P������� ��?�ί�u����(� ��Ͽ^�󿂿�)ϸ� M�ܿqσ�ϧ�6��� Z�l�ߐ�%ߴ��[� ���ߣߵ�D���h� ����3���W����� ����@����v�� ��/�A���e������ *���N���r����� =��6s�&� �\��'�K �o��4�X ���#/�G/Y/� }//�/�/B/�/f/�/ �/�/1?�/U?�/N?�? ?�?>?�?�?t?	O�? -O?O�?cO�?�OO(O��O�F�$FILE�_DGBCK 1�]���@��� < ��)
SUMMAR�Y.DG�OsLM�D:�O;_@D�iag Summ�ary<_IJ
CONSLOG1__&Q�_�_NQConsole log�_�HK	TPACCNĵ_o%o?oJUT�P Accoun�tin�_IJFR�6:IPKDMPO.ZIPsowH
�o��oKU[`Excep�tion�oyk'PMEMCHECK5o�_*_K�QMem�ory Data|L�F1l�)6qRIPE�_$6��Zs%�q Pa?cket L�_�D�L�$�	r�qST�AT���S� �%�rStat�usT��	FTP����:���Vw�Qm�ment TBD�؏� >I)E?THERNE����
q�[�NQEth�ern�p�Pfig�ura�oODDCSVRF̏��ďݟ�d��� veri?fy all��{D��.���DIFF�՟��͟b��s��di�ffd��
q��CHG01Y�@�R��f�Xz���-?��2ݯ�į֯k�v�����3pa�H�Z�� ���ϥ�VTRND?IAG.LS�̿�޿s�^q3� Op�e���q SQnos�ticEW��)�VDEV7�DA�Tt�Q�c�u�g�V�is��Devic9e�Ϫ�IMG7ºo�����y��s�Imsagߨ�UP���ES��T�FRS�:\�� �OQUp�dates Li�st �IJg�FL?EXEVENQ�X��j߃�f�F� UI�F Ev���B,��s�)
PSRBWLD.CM���sL������PPS�_ROBOWEL���GLo�GRAP?HICS4Dy�b��t��%4D �Graphics� Fileu��AOwɿ�rGIG����u�
YvGig�E�ة�BN�? �)��HADOW������\sSh�adow Chasng���vbQ?RCMERR�n�\s� CFG� Error�t�ail� MA���CMSGLIB��"^o�� ��T�)�ZD����/Xw7ZD6 ad�H=PNOTI����
/�/ZuNoti�fic��H/��AGUO�/yO?�O'?P? OOt??�?�?9?�?]? �?O�?(O�?LO^O�? �OO�O5O�O�OkO _ �O$_6_�OZ_�O~_�_ _�_C_�_�_y_o�_ 2o�_?oho�_�oo�o �oQo�ouo
�o@ �odv�)�M �����<�N�� r������7�̏[��� ���&���J�ُW��� ���3�ȟڟi����� "�4�ßX��|���� ��A�֯e�����0� ��T�f���������� O��s��ϩ�>�Ϳ b��oϘ�'ϼ�K��� �ρ�ߥ�:�L���p� �ϔߦ�5���Y���}� ��$��H���l�~�� ��1�����g���� � 2���V���z�	����� ?���c���
��.�� Rd�����M �q�<�` ���%�I�� /�8/J/�n/� �/!/�/�/W/�/{/? "?�/F?�/j?|??�?�/?�?�?�$FIL�E_FRSPRT�  ���0�����8M�DONLY 1]��5�0 
 ��)MD:_VD�AEXTP.ZZ�Z�?�?_OnK6�%NO Back file 9O�4S�6Pe?�OOO �O�?�O__?>_�Ob_ t__�_'_�_�_]_�_ �_o(o�_Lo�_po�_ }o�o5o�oYo�o �o $�oHZ�o~� �C�g��	�2� �V��z������?� ԏ�u�
���.�@��4?VISBCKHA>&C*.VDA������FR:\Z�I�ON\DATA\�v����Vis?ion VD�B�� ŏ���'�5��Y�� j������B�ׯ�x� ���1���үg����� ��X���P��t���� ��?�οc�u�ϙ�(� ��L�^��ς��)��� M���q� ߂ߧ�6��� Z�����%��I��������:LUI_C�ONFIG ^��5m��� $ h�F{�5�������)�;�I���|x q�s�����������a� �� $6��Gl ~���K���  2�Vhz� ��G���
// ./�R/d/v/�/�/�/ C/�/�/�/??*?�/ N?`?r?�?�?�???�? �?�?OO&O�?JO\O nO�O�O)O�O�O�O�O �O_�O4_F_X_j_|_ �_%_�_�_�_�_�_o �_0oBoTofoxo�o!o �o�o�o�o�o�o, >Pbt��� �����(�:�L� ^�p��������ʏ܏ ���$�6�H�Z�l� �������Ɵ؟ꟁ� � �2�D�V�h����� ����¯ԯ�}�
�� .�@�R�d��������� ��п�y���*�<� N�`����ϖϨϺ��� ��u���&�8�J��� [߀ߒߤ߶���_��� ���"�4�F���j�|� ������[������ �0�B���f�x����� ����W�����, >��bt���� O��(:��  xFS��$FLUI_DA�TA _��}����uRESULT �2`�� ��T�/wiz�ard/guid�ed/steps/Expertb ��//+/=/O/a/�s/�/�/�*�Co�ntinue w�ith G�ance�/�/�/??(?�:?L?^?p?�?�?�? �T-U��90 �� �?���9��ps�?0OBO TOfOxO�O�O�O�O�O �O�O� �_/_A_S_ e_w_�_�_�_�_�_�_@�_n�?�?�?�<Frip�Oo�o�o �o�o�o�o�o!3 E_i{���� �����/�A�S� o$on�HoAO��TimeUS/DST[������+��=�O�a�s������'Enabl�/˟ݟ ���%�7�I�[�m�(�����T�?{�0ݯ����Æ24Ώ3� E�W�i�{�������ÿ տ翦����/�A�S� e�wωϛϭϿ����� �ϴ�Ưد� G��?Region�χ� �߽߫����������)�;�+Americasou���� ����������)�;��?�y�#߅�G�Y�>�ditorL��� ����#5GYk�}��+ Touc�h Panel ��� (recommen�)��� *<N`r��U��e�w������>��accesd�./ @/R/d/v/�/�/�/�/��/�/Q|Conn�ect to N?etwork�/(? :?L?^?p?�?�?�?�?P�?�?�?Y���������!/��Introducts� �O�O�O�O�O�O�O_ _(_:_U^_p_�_�_ �_�_�_�_�_ oo$o6oHo e�Oeo?O �X_�o�o�o�o '9K]o��R_ ������#�5�@G�Y�k�}�����h`�ooj}oߏ�o�� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ쯫���Ϗ1��X� j�|�������Ŀֿ� ����0��A�f�x� �ϜϮ���������� �,�>���_�!���E� �߼���������(� :�L�^�p���߸� ������ ��$�6�H� Z�l�~���O߱�s��� ���� 2DVh z�������� 
.@Rdv� �������/�� '/���`/r/�/�/�/ �/�/�/�/??&?8? �\?n?�?�?�?�?�? �?�?�?O"O4O�UO /yO�OO?�O�O�O�O �O__0_B_T_f_x_ �_I?�_�_�_�_�_o o,o>oPoboto�oEO �OiO�o�o�O( :L^p���� ���_ ��$�6�H� Z�l�~�������Ə؏ �o�o�o�/��oV�h� z�������ԟ��� 
��.��R�d�v��� ������Я����� *��������C��� ��̿޿���&�8� J�\�nπ�?��϶��� �������"�4�F�X� j�|ߎ�M�_�q��ߕ� ����0�B�T�f�x� ������������ �,�>�P�b�t����� ���������߱���% ��L^p���� ��� $��5 Zl~����� ��/ /2/��S/ w/9�/�/�/�/�/�/ 
??.?@?R?d?v?�? �/�?�?�?�?�?OO *O<ONO`OrO�OC/�O g/�O�/�O__&_8_ J_\_n_�_�_�_�_�_ �_�?�_o"o4oFoXo jo|o�o�o�o�o�o�O �o�O�O�oTfx �������� �,��_P�b�t����� ����Ώ�����(� �oI�m��C����� ʟܟ� ��$�6�H� Z�l�~�=�����Ưد ���� �2�D�V�h� z�9���]���ѿ���� 
��.�@�R�d�vψ� �ϬϾ��Ϗ����� *�<�N�`�r߄ߖߨ� ���ߋ�տ����#�� J�\�n������� �������"���F�X� j�|������������� ��������u 7������ ,>Pbt3�� �����//(/ :/L/^/p/�/ASe �/��/ ??$?6?H? Z?l?~?�?�?�?�?� �?�?O O2ODOVOhO zO�O�O�O�O�O�/�/ �/_�/@_R_d_v_�_ �_�_�_�_�_�_oo �?)oNo`oro�o�o�o �o�o�o�o&�O G	_k-_���� ����"�4�F�X� j�|������ď֏� ����0�B�T�f�x� 7��[������ �,�>�P�b�t����� ����ί�����(� :�L�^�p��������� ʿ��뿭��џӿH� Z�l�~ϐϢϴ����� ����� �߯D�V�h� zߌߞ߰��������� 
��ۿ=���a�s�7� ������������ *�<�N�`�r�1ߖ��� ��������&8 J\n-�w�Q�� ����"4FX j|������� �//0/B/T/f/x/ �/�/�/�/���/ ?�>?P?b?t?�?�? �?�?�?�?�?OO� :OLO^OpO�O�O�O�O �O�O�O __�/�/�/ ?i_+?�_�_�_�_�_ �_�_o o2oDoVoho 'O�o�o�o�o�o�o�o 
.@Rdv5_ G_Y_�}_���� *�<�N�`�r������� ��yoޏ����&�8� J�\�n���������ȟ �����4�F�X� j�|�������į֯� ���ˏ�B�T�f�x� ��������ҿ���� �ٟ;���_�!��Ϙ� �ϼ���������(� :�L�^�p߁ϔߦ߸� ������ ��$�6�H� Z�l�+ύ�Oϱ�s��� ����� �2�D�V�h� z��������������� 
.@Rdv� ���}������ �<N`r��� ����//��8/ J/\/n/�/�/�/�/�/ �/�/�/?�1?�U? g?+/�?�?�?�?�?�? �?OO0OBOTOfO%/ �O�O�O�O�O�O�O_ _,_>_P_b_!?k?E? �_�_{?�_�_oo(o :oLo^opo�o�o�o�o wO�o�o $6H Zl~���s_�_ �_���_2�D�V�h� z�������ԏ��� 
��o.�@�R�d�v��� ������П����� ���]�������� ��̯ޯ���&�8� J�\����������ȿ ڿ����"�4�F�X� j�)�;�M���q����� ����0�B�T�f�x� �ߜ߮�m�������� �,�>�P�b�t��� ���{ύϟ����(� :�L�^�p��������� ������ ��6H Zl~����� ����/��S� z������� 
//./@/R/d/u�/ �/�/�/�/�/�/?? *?<?N?`?�?C�? g�?�?�?OO&O8O JO\OnO�O�O�O�Ou/ �O�O�O_"_4_F_X_ j_|_�_�_�_q?�_�? �_�?�_0oBoTofoxo �o�o�o�o�o�o�o �O,>Pbt�� �������_%� �_I�[��������� ʏ܏� ��$�6�H� Z�~�������Ɵ؟ ���� �2�D�V�� _�9�����o�ԯ��� 
��.�@�R�d�v��� ����k�п����� *�<�N�`�rτϖϨ� g�����������&�8� J�\�n߀ߒߤ߶��� �����߽�"�4�F�X� j�|���������� ���������Q��x� �������������� ,>P�t�� �����( :L^�/�A��e� ��� //$/6/H/ Z/l/~/�/�/a�/�/ �/�/? ?2?D?V?h? z?�?�?�?o���? �O.O@OROdOvO�O �O�O�O�O�O�O�/_ *_<_N_`_r_�_�_�_ �_�_�_�_o�?#o�? Go	Ono�o�o�o�o�o �o�o�o"4FX io|������ ���0�B�T�ou� 7o��[o��ҏ���� �,�>�P�b�t����� ��iΟ�����(� :�L�^�p�������e� ǯ��믭���$�6�H� Z�l�~�������ƿؿ ����� �2�D�V�h� zόϞϰ��������� ���ۯ=�O��v߈� �߬߾��������� *�<�N��r���� ����������&�8� J�	�S�-�w���c��� ������"4FX j|��_���� �0BTfx ��[�������� /,/>/P/b/t/�/�/ �/�/�/�/�/�?(? :?L?^?p?�?�?�?�? �?�?�?����EO /lO~O�O�O�O�O�O �O�O_ _2_D_?h_ z_�_�_�_�_�_�_�_ 
oo.o@oRoO#O5O �oYO�o�o�o�o *<N`r��U_ ������&�8� J�\�n�������couo �o鏫o�"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү����� �ُ;���b�t����� ����ο����(� :�L�]�pςϔϦϸ� ������ ��$�6�H� �i�+���O������� ����� �2�D�V�h� z���]��������� 
��.�@�R�d�v��� ��Y߻�}����ߣ� *<N`r��� ������&8 J\n����� ����/��1/C/ j/|/�/�/�/�/�/�/ �/??0?B?f?x? �?�?�?�?�?�?�?O O,O>O�G/!/kO�O W/�O�O�O�O__(_ :_L_^_p_�_�_S?�_ �_�_�_ oo$o6oHo Zolo~o�oOO�OsO�o �o�O 2DVh z�������_ 
��.�@�R�d�v��� ������Џ⏡o�o�o �o9��o`�r������� ��̟ޟ���&�8� �\�n���������ȯ گ����"�4�F�� �)���M���Ŀֿ� ����0�B�T�f�x� ��I������������ �,�>�P�b�t߆ߘ� W�i�{��ߟ���(� :�L�^�p����� ��������$�6�H� Z�l�~����������� ������/��Vh z������� 
.@Qdv� ������// */</��]/�/C�/ �/�/�/�/??&?8? J?\?n?�?�?Q�?�? �?�?�?O"O4OFOXO jO|O�OM/�Oq/�O�/ �O__0_B_T_f_x_ �_�_�_�_�_�_�?o o,o>oPoboto�o�o �o�o�o�o�O�O% 7�_^p���� ��� ��$�6��_ Z�l�~�������Ə؏ ���� �2��o; _���K��ԟ��� 
��.�@�R�d�v��� G�����Я����� *�<�N�`�r���C��� g���ۿ����&�8� J�\�nπϒϤ϶��� �ϙ����"�4�F�X� j�|ߎߠ߲����ߕ� ����˿-��T�f�x� ������������� �,���P�b�t����� ����������( :����A�� ��� $6H Zl~=����� ��/ /2/D/V/h/ z/�/K]o�/��/ 
??.?@?R?d?v?�? �?�?�?�?��?OO *O<ONO`OrO�O�O�O �O�O�O�/�O�/#_�/ J_\_n_�_�_�_�_�_ �_�_�_o"o4oE_Xo jo|o�o�o�o�o�o�o �o0�OQ_u 7_������� �,�>�P�b�t���Eo ����Ώ�����(� :�L�^�p���A��e ǟ��� ��$�6�H� Z�l�~�������Ưد ����� �2�D�V�h� z�������¿Կ���� ���+��R�d�vψ� �ϬϾ��������� *��N�`�r߄ߖߨ� ����������&�� /�	�S�}�?Ϥ���� �������"�4�F�X� j�|�;ߠ��������� ��0BTfx 7��[����� ,>Pbt�� ������//(/ :/L/^/p/�/�/�/�/ �/����!?�H? Z?l?~?�?�?�?�?�? �?�?O O�DOVOhO zO�O�O�O�O�O�O�O 
__._�/�/?s_5? �_�_�_�_�_�_oo *o<oNo`oro1O�o�o �o�o�o�o&8 J\n�?_Q_c_� �_���"�4�F�X� j�|�������ď�oՏ ����0�B�T�f�x� ��������ҟ�� ��>�P�b�t����� ����ί����(� 9�L�^�p��������� ʿܿ� ��$��E� �i�+��Ϣϴ����� ����� �2�D�V�h� z�9��߰��������� 
��.�@�R�d�v�5� ��Yϻ�}������ *�<�N�`�r������� ��������&8 J\n����� �������FX j|������ �//��B/T/f/x/ �/�/�/�/�/�/�/? ?�#�G?q?3�? �?�?�?�?�?OO(O :OLO^OpO//�O�O�O �O�O�O __$_6_H_ Z_l_+?u?O?�_�_�? �_�_o o2oDoVoho zo�o�o�o�o�O�o�o 
.@Rdv� ���}_�_�_�_� �_<�N�`�r������� ��̏ޏ�����o8� J�\�n���������ȟ ڟ����"���� g�)�������į֯� ����0�B�T�f�%� ��������ҿ���� �,�>�P�b�t�3�E� W���{�������(� :�L�^�p߂ߔߦ߸� w����� ��$�6�H� Z�l�~������� ������2�D�V�h� z��������������� 
-�@Rdv� ������ ��9��]���� ����//&/8/ J/\/n/-�/�/�/�/ �/�/�/?"?4?F?X? j?)�?M�?qs?�? �?OO0OBOTOfOxO �O�O�O�O/�O�O_ _,_>_P_b_t_�_�_ �_�_{?�_�?oo�O :oLo^opo�o�o�o�o �o�o�o �O6H Zl~����� ����_o�_;�e� 'o������ԏ��� 
��.�@�R�d�#�� ������П����� *�<�N�`��i�C��� ��y�ޯ���&�8� J�\�n���������u� ڿ����"�4�F�X� j�|ώϠϲ�q����� ��	�˯0�B�T�f�x� �ߜ߮���������� ǿ,�>�P�b�t��� ������������� ����[�߂������� ������ $6H Z�~����� �� 2DVh '�9�K��o���� 
//./@/R/d/v/�/ �/�/k�/�/�/?? *?<?N?`?r?�?�?�? �?y�?��?�&O8O JO\OnO�O�O�O�O�O �O�O�O_!O4_F_X_ j_|_�_�_�_�_�_�_ �_o�?-o�?QoOxo �o�o�o�o�o�o�o ,>Pb!_�� �������(� :�L�^�o�Ao��eo g�܏� ��$�6�H� Z�l�~�������s؟ ���� �2�D�V�h� z�������o�ѯ���� �˟.�@�R�d�v��� ������п����ş *�<�N�`�rτϖϨ� ������������� /�Y���ߒߤ߶��� �������"�4�F�X� �|���������� ����0�B�T��]� 7߁���m������� ,>Pbt�� �i����( :L^p���e� w��������$/6/H/ Z/l/~/�/�/�/�/�/ �/�/� ?2?D?V?h? z?�?�?�?�?�?�?�? 
O���OO/vO�O �O�O�O�O�O�O__ *_<_N_?r_�_�_�_ �_�_�_�_oo&o8o Jo\oO-O?O�ocO�o �o�o�o"4FX j|��__��� ���0�B�T�f�x� ������moϏ�o�o �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ���!��E� �l�~�������ƿؿ ���� �2�D�V�� zόϞϰ��������� 
��.�@�R��s�5� ��Y�[��������� *�<�N�`�r���� g���������&�8� J�\�n�������c��� ��������"4FX j|������ ���0BTfx ��������� ����#/M/t/�/�/ �/�/�/�/�/??(? :?L?p?�?�?�?�? �?�?�? OO$O6OHO /Q/+/uO�Oa/�O�O �O�O_ _2_D_V_h_ z_�_�_]?�_�_�_�_ 
oo.o@oRodovo�o �oYOkO}O�O�o�O *<N`r��� �����_�&�8� J�\�n���������ȏ ڏ����o�o�oC� j�|�������ğ֟� ����0�B��f�x� ��������ү���� �,�>�P��!�3�������$FMR2_�GRP 1a���� ��C4  B�[�	� [�߿�ܰE�� F@ �ǂ5W�S�ܰJ���NJk�I'�PKHu��IP��sF!���?ǀ  W�S�ܰ9��<9�8�96C'6<�,5���Ag�  �Ϲ�BHٳ�B�հ����@�3]3�33S�۴x��ܰ@UUT'��@��8��W�>u.��>*��<�����=[�B=����=|	<��K�<�q�=��mo���8��x	7H<8��^6�Hc7��x?�����������"��F�X���_CF�G b»T �Q����X�NO� º
F0��� ��W�RM_C�HKTYP  ���[�ʰ̰����RO=M�_MIN�[�W��9����X���SSBh�c�� ݶf�[��]����^�TP_D�EF_O�[�|ʳ��IRCOM�����$GENOV_RD_DO.�d�n��THR.� d�d��_ENB�� ���RAVC��d�O�Z� ���F�s  G!� G�Ƀ�I�C�I(i J���+��%����� [�QOU��j¼�������<6�i�C�;]�~[�C�  D��+��@���B�����.��R SMT��k_	ΰ\��$HOSTCh�s1l¹[��d��۰ MC[����/Z�  27�.0� 1�/  e�/??'?9?G:�/�j?|?�?�?�,Z?T3	�anonymou y �?�?	OO-O?N�/ڰRHRK�/�?�O�/ �O�O�O�O_V?3_E_ W_i_�O&_�?�_�_�_ �_�_@O�_dOvOSo�_ �Ojo�o�o�o�o_�o +=`o�_�_� ����o&o8oJo L9��o]�o������� �oɏۏ����4�j +�Y�k�}������� �� ��T�1�C�U� g�����������ӯ�� x�>��-�?�Q�c��� ��Ο���Ͽ��� �)�;ς�_�qσϕ� ��ʿ ������%� 7�~�����߶ϣ�� ���������Ϻ�3�E� W�i�ߍ��ϱ����� ����@�R�d�v�x�J� �߉������������ +=`���������:$h!EN�T 1m P�!V  7  ?.c&�J� n���/�)/� M//q/4/�/X/j/�/ �/�/�/?�/7?�/? m?0?�?T?�?x?�?�? �?O�?3O�?WOO{O >O�ObO�O�O�O�O�O _�OA__e_(_:_�_�^_�_�_�_�ZQUICC0�_�_�_?o�d1@oo.o�od2�olo~o�o!ROUTER�o�o�o/!PCJOG0�!192.�168.0.10�	o�SCAMPRT,�\!pu1yp���vRT�o��� �!Softwa�re Opera�tor Pane�l�mn��NAM�E !�
!R�OBO�v�S_C�FG 1l�	 ��Aut�o-starte�d'�FTP2� �I�K2��V�h�z� ������ԟ���� 	���@�R�d�v���	� ������:���)� ;�M�_�&��������� ˿�p���%�7�I� [��"�4�F�ڿ��� �����!�3���W�i� {ߍߟ���D������� ��/�vψϚ�w�� ���Ͽ��������� +�=�O�a�������� ��������8�J�\�n� p�]������ ����#5X� k}���� 0/D1/xU/g/y/ �/RH/�/�/�/�// ?�/??Q?c?u?�?� ��/?�?:/O)O ;OMO_O&?�O�O�O�O �O�?pO__%_7_I_ [_�?�?�?t_�O�_O �_�_o!o3o�OWoio {o�o�_�oDo�o�o�o�����_ERR� n��-=vPDUSIZ  �`�^�P�Tt>muW�RD ?΅�Q��  guest�f�������~�SCDMN�GRP 2o΅;Wp��Q�`����fKL� 	P01.05 8�Q�   �|���  ;|�� � z[ ����w���*���}Ť�x����`[ݏȏ��בP�Ԡ������)�����D�r���U؊p"�Pl�P���	Dx��dx�*������%�_GROU7�p*LyN��	/�o�.��QUP��UTuY� �TYàL}�?pTTP_AU�TH 1qL{ �<!iPend�an����o֢!�KAREL:*8������KC��ɯ�ۯ��VISION SET�9�� ��P�>�h��f�����������ҿ�����X�CTRL r�L}O�uſa
��kFFF9E3-���TFRS:DE�FAULT���FANUC We�b Server �ʅ�t�X���t@����1�C�U�g�;tWR�_CONFIG ;s;� ��=q�IDL_CPU_kPC���aBȠP��� BH��MIN��܅q��GNR_I�OFq{r�`Rx��NP�T_SIM_DO���STAL_oSCRN� �.��INTPMODN�TOLQ����RT�Y0����-�\�EN�BQ�-���OLN/K 1tL{�p������)�;�M���M�ASTE�%���SLAVE uL�|�RAMCACH�Ek�c�O^�O_CcFG������UOC������CMT_OPp���PzYCL�������_ASG 19v;��q
 O�r ��������&8J\W�EN�UMzsPy
��I�P����RTRY_CN��M�=�zs����Tu ������w����p/�p��P_M�EMBERS 2Yx;�l� $��X"���?�Q'W/i)��R�CA_ACC 2�y�  X�c�� ˣ t�� /�` 5!�@�`���`�&4��C�6��/�$  ��b�,�$BUF0�01 2z�= �`�u0  uW0`�:4�:4�:4��:3aZ4Z4-�Z4=Z4NZ4`Z4p�Z4�Z4�Z4�Z4��Z4�Z4�Z4�Z4�V:3b�4�4+�4U:�4L�4\�4n�4��x�xbQ4b��:3c"D"D/�"DA"DR"Dd"Dt*"D�"D�"D�"D94�cA4c�b�  �b�^2u0:1^~I@k�	x^r�D�h�h�@^�L�hLh  _2K�xK@_rkXc���` Y�@YW�`:4!:41:4�B:4ID`QD`YD`�aD`�:4�:392 $?63:1@1ERI0ERQ0 ERY0:1`1eRi0eRq0 eRy0eR�0eR�0eR�0 eR�0eR�0eR�0eR�0 eR�0eR�0eR�0eR�0 :1�1�R�0�R�0�R�0 �R�0�R@�R	@�R@<AAY�x A:1 (A-b1@-b9@-bA@-b I@-bQ@-bY@-ba@-b i@-bq@-bBT�A-b�@`�A�I�B�O�NkXGP �@�A�AER�@ER�@ER �@ERRd�AERbdQER PERP:193-_65 GSNrI2WSNrY2gSnr i2wSnry2�Snr�2�S nr�2�Snr�2�Snr�2 �Snr�2�S���3�S�r �2�S�r�2c�r	Bc �rct C/c6�1B?c6� ABOc6�QB_c6�aBoc 6�qBc6�St�C�c�� [��a���`���`���A Ƃ�@Nr�B�cNr�B�c Nr�B�cNrc� SsNr`Rs�Ԝ!��2{�Q4r�}ŋ���<��௑o�o��2�HIS�!2}� ܷ!� 2024-07-2O�����П�v��  8�;  Ղ:�`��" *�!N����+�=�O�a�o�X�b꩘2������Ư0د���m�b�l��p�)�;�r��fn��6-27��~���������fn�������"�}��ga�6 m�Z�l�~ϵ�o�Ղo�ѵgۿ��������.}��j�a�5I�6��H�Zߵ� 7 ɽł�j���߲߸����y��cNa�1ട�#�5�� 9� ��cN�߀���\��}��mva�0H�`��������Z�M g9 �@D�mvL�;M Y�k�}���r�� ,P����������'�%,r�J�`r�c�9
� :��d_q� q���������;L�b��o�M:L ^�^�����(�96d>dٰ%/ $/6/H/6���~/�/�/ $�"�`"���/�/  ??$?�$�Z?l?~?��:��@��� ��?�?�?�?����O@COUOgO. �2�2�P �m��?�O�O�O�O���m/_$_6_$�& # @�A�c�2Q�o�cD_�_�_�_�� 3r����_o$o6o'��Td��ecro �o�o�o��o�o&�&�AsN` r�r��o��� )�Br� Br?uٰJ7� I�[�m�[/_����Ǐ ����&��%�7�I�@7?I?�����$�Wd ƒƒnPBr����� 	��	OOv�c�u����,�Wd��gbN ����Я����O�OO��<�N�`�)�Xc(�A�ה��Q�i���¿Կ��__I_CFG �2~�[ H
�Cycle Ti�me(�Bus}y�Idl�^-�min�S��Up� �R�ead(�DoqwG�C�W���Count �	N'um �.������(�����PROG����U�P��)/softpa�rt/genli�nk?curre�nt=menup�age,1133,1�C�U�g�y�T����SDT_ISO�LC  �Y� ����J23_D�SP_ENB  ���V���INC ����(���A  � ?�  =�̟�<#�
���:�o �2�D�(�X/�l���OB��C���O��ֆ�G_GR�OUP 1���}�"< ���P����t�?����(�Q'�L�^�p�/� ���������\�~��G_IN_AUT�O����POSRE����KANJI_�MASK0��DR�ELMON ��[��(�y���������f�Ã�����(�-��KCwL_L NUM���G$KEYLOGOGINGD�P�������LANGUA_GE �U���DEFAUgLT ��QLG������S��(�x�ఔ�8T�H  -�(�'0縤(��1x��K�(�;��
*!(UT1:\ J/ L/Y/k/}/�/��/�/�/�/�/�/$>(��H?�VLN_DISP ���P�&�|$�^4OCTOLĔ�Dz����
�1GB?OOK ���A 1V�11�@��% O!O3OEOWOiKyM�TËIgF	�5)������O}���2_BU�FF 2��� ��[�e_�2�� 6_M�R_d_�_�_�_�_ �_�_�_�_o3o*o<o No`o�o�o�o�o���A?DCS ����� �L�O��+=O|a�dIO 2��k� ������ �������� *�:�L�^�r������� ��ʏ܏���$�6��J�uuER_ITM��d������ǟٟ� ���!�3�E�W�i�{� ������ïկ������7x�SEVD��.t�TYP����s�p�����)RSTe��eSCRN_FLW 2��}��� ��/�A�S�e�wϨ��TP{��b��=NGNAM��E��d7UPSf0GI��2�����_LOA�D��G %��%�DROP_�E�ITO_3�ϑ�MAXUALRMb,2�@���
K���'_PR��2  �3�AK�Ci0��qO=_x'X�Ӭ�P 2��;W �*V	����
* ���4��*� �'�`�	xN��z�� ����������1�C� &�g�R���n������� ����	��?*c FX������ �;0q\ �������/ �/I/4/m/X/�/�/ �/�/�/�/�/�/!?? E?0?i?{?^?�?�?�? �?�?�?�?OOAOSO�6OwObO�OD�DBG*� ��գѢѤO��@_LDXDIS�A����ssMEMO�_AP��E ?��
 �Ax$_ 6_H_Z_l_~_�_�_K��FRQ_CFG k����CA w�@��S�@<��d%��\o�_�P�Ґ��{��*Z`=/\b **:eb�D Xojho�F�o�o�o�o �o�o;�O��d�Z�U�y|��z,( 9�Mt���1�� B�g�N���r���������̏	���?�A�I�SC 1���K` ��O�����O���O֟�����K�]�_MST�R �3��SC/D 1�]��l� �{�����دïկ ���2��V�A�z�e� ������Կ������ �@�+�=�v�aϚυ� �ϩ���������<� '�`�K߄�oߨߓߥ� �������&��J�5� Z��k�������� ������F�1�j�U� ��y��������������0T?x�M�K�Q�,��Q�$�MLTARM�Ru�?g� ~s��@���@METP�U�@l��4�N�DSP_ADCO�L�@!CMNT�7(FNSWiS7TLIx *%� �,����Q�|�*POSCF�=�PRPMV��ST51�,� 4�R#�
g!|qg% w/�'c/�/�/�/�/�/ �/?�/?G?)?;?}? _?q?�?�?�?�?�1*�SING_CHK�  {$MODA�S�e���#E�DEV 	�J	�MC:WLHSI�ZE�Ml �#ETA�SK %�J%$�12345678�9 �O�E!GTRI�G 1�,� l �Eo#_�y_S_�}�F�YP�A�u9D"CE�M_INF 1��?k`)AT?&FV0E0X_�]�)�QE0V1&�A3&B1&D2�&S0&C1S0}=�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_�_o �3o��o���o� �"�4��X��� ASe֏���C� 0���f�!���q��� ��s�䟗�����͏>� �b���s���K���w� ��ٯ�ɟ۟L��� �#�����Y�ʿ�� ����$�߿H�/�l�~� 1���U�g�y����ϯ�  �2�i�V�	�z�5ߋ��ߗ���PONITO�R�G ?kK  � 	EXEC�1o�2�3�4��5��@�7�8
�9o��� ��(��4��@��L� ��X��d��p��|⪂�2��2��2��2���2��2��2��2���2��2��3��3��3(�#AR_GRP_SV 1��[� (�1?�}��*�����@(�������,&�RM�A_D�sҔN��ION_D�B-@�1Ml  �l ]FH"- -	��l FH��N �BL"FI-ud�1}E���)PL�_NAME !��E� �!De�fault Pe�rsonalit�y (from �FD)b*RR2��� 1�L�X�L�p�X  d�-?Qcu �������/ /)/;/M/_/q/�/�/�/f2)�/�/�/?�?,?>?P?b?t?f< �/�?�?�?�?�?�?
O�O.O@OROdOc	�6D�?�N
�O�OfP�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ �O�O2oDoVohozo�o �o�o�o�o�o�o
 .@o!ov��� ������*�<��N�`�r����� �Fs  GT��G�Me��x �ÏՍfd������ �(�6������
 �m�p~�h����� �� ����ğ֟�����:����
�]�m�f��	�`������į��:�oAb	����� A�  /� ��P����r������� ^�˿ݿȿ��%���R�� 1��	X ���, � ���� a� @D� M t�?�z�`�?f <|�fA/��t�{	ު�;�	l��	 ��x�J���� � �� ��<�@���� ���·�K�K� ��K=*�J����J���J9��
�ԏC����@�t�@{S�\��(Ehє���.��I���}ڌ���T;f�����$��3��´7  �@��>�Թ��$�  >�����ӧUf��x`���� �
����Ǌ��� �  �{  @T������  �H ��l�ϊ�-�	'� �� ��I� ?�  �<�+��:�È��È=G�����0Ӂ��N ��[��n @@���f���f�k����,�av�  '���Yэ�@2��@��0@�Ш����C��Cb C��\�C������G�K@������� )�Bb $/�!��L��Dz�o�ߓ~���0��( ?�� -���`������!���/�����恀?�fafG�*<� }��q�1�8����>���bp��(�(���P���	������>�?�����x���W�<�
6b<߈;�܍�<�ê<���<�^��dI/��A�{��f�|��,�?fff?_��?&� T�@�.��"�J<?�\��"N\�5���!�� (�|��/z��/j'��[ 0??T???x?c?�?�?��?�?�?�?5��%F ��?2O�?VO�/wO�)�IO�OEHG@ G�@0��G�� G}ଙO�O�O_	_B_�-_f_Q_BL��B��Aw_[_�_b��_�[ �_��mO3o�OZo�_~o�o�o�o���b��PV( @|po	lo@-*cU�ߡA���r5eCP�Lo�}?����#�l�5��W�s��6�3Cv�q�CH3� jD�t����q�����|^�(hA� �A�LffA]��??�$�?��;��°u�æ�)��	ff��Cϼ#�
���g\�)�"�33C�
������<����؎G�B����L�B�s����	"�;�H�ۚG���!G��WIY�E���C�+��8�I۪I��5�HgMG��3E��RC��j=x�
�pI����G��fIV�=�E<YD �C<�ݟȟ����7� "�[�F��j������� ٯį���!��E�0� i�T�f�����ÿ��� ҿ����A�,�e�P� ��tϭϘ��ϼ���� ��+��O�:�s�^߃� �ߔ��߸������ � 9�$�6�o�Z��~�� �����������5� � Y�D�}�h����������������
C.(�䁳��/"��<�<��t��q3�8����q�4Mgu���q��VwQ�
4p�+4�]$$d@R�v���uPD"	P��Q�_/Z/0=/(/a/L+Rg/n/`�/�/�/�/�/  %��/�/+??O?:?s?�/�_�?�?�?�; �?�?O�? OFO4O�rLO^O�O�O�O�O�O��J  2 FsޖwGT�V��M�uBO�|r�pp�C��S@�R_�poy_��_^_�_o \!�WɃ�_oo(o~�z?���@@�z��D�p�pk1:�p�~
 6o�o �o�o�o�o�o)�;M_q�ڊsa �����D���$MR_CABL�E 2�� S]��T�La�Ma?�PMaLb�p��Z��&P�C�p�!O4>�B����"כ��� >�!F�?��F��"�~�v�l  ��&Py�v�wdN�{0���$ �� z�RefF�[(�7�I�XT��6P� ;C$�Č�$���Q� F�?U	F.�,���|% ��&P��C����=�������Q�S�	F�hڅ��s9�"T�p� �J�D�V�h�z�ߟڟ ����ԟ�K�
��F��@�R�d��	j��#�  ������;h�H�Z��l�;h*��**} �sOM ��y����� j �l�%% 23�45678901�ɿ۵ ƿ���� ��� AQ� �!
��z�not s�ent ���W��TESTF�ECSALG� e�g�ZAQd��ga%�
,���@���$�r�̹������� 9�UD1:\mai�ntenance�s.xmS�.�@��vj�DEFA�ULT�\�rGRP� 2���  p�� �J�%  �%�1st mec�hanical �check��!����������E ��Z�(�:�L�^��"���controller�Ԍ��߰��D����� ��$�s�cM��L��""8b���v��B�����������/�C}�a�6����dv����s�C��ge��.� battery�&��E	S(:�L^p�	|�dui�z�ablet  �D�а�R������/"/4/s�>�greas��'f�r#-� |!�/�E��/�/�/�/�/s�
�oi,�g/y/�/�/t?�?�?�?�?"s��
�XֈW��1!<X�AO�E
c?8O JO\OnO�O�t��?O��'O�O_ _2_�D_s�Overh�auE��L��R !xXЌQ�_���O�_ �_�_�_oX�$�_0o ϤFi4oVٰ_�o�o�o �o�oo�o@oRodo% K]o���o� *��#�5�G�� X�}�����ŏ׏� ���\�1�C���g��� ��������ӟ"���F� X�-�|�Q�c�u����� 蟽����B��)� ;�M�_�����ү䯹� �ݿ���%�t�I� �����ο�ϵ����� ��:��^�pςϔ�i� {ߍߟ߱� ���$�6� H�	�/�A�S�e�w��� ������������� +�z�<�a���d���� ��������@�'v� K��o���� �*<`5GY k}����& �//1/C/�g/� ��/��/�/�/�/	? X/-?|/�/c?�/�?�? �?�?�??�?B?T?f? x?MO_OqO�O�O�?�O OO,O�O_%_7_I_ [_�O_�O�O�O�_�_��_�_o!o�T	 T "oOoaoso�_�o�_�k �o�o�o�o�o�o2D z��`r� ����.�@��� v�����\�n�Џ⏤�����R ��Q?�  @�a  �oW�i�{��fC������̟aX*�**  ������ �2�D���h�z������� �_�S������կ 7�I�[�����ɯ/��� ǿٿ#���!�3�}� ����{ύϟ��s��� ����C�U�g��S�e� w�9ߛ߭߿�	�߉e��a�$MR_H�IST 2������ 
 \jR$� 2345678�901*�2����)�9c_���R��a_ ���������=�O�a� �*�x�����r����� ��9��]o& �J����� #�G�k}4���d�SKCFMA�P  ��R�����`���ONREL  �����лE�XCFENB'
8��!FNC$/$�JOGOVLIM�'d�m �KEY�'p%y%_PA�N(�"�"�RUN�`,�+SFSPD�TYPD(%�SI�GN/$T1MO�Tb/!�_CE_GRP 1����"�:`��n?�c [?�?�؆?�?~?�?�? �?!O�?EO�?:O{O2O �O�OhO�O�O�O_�O /_�O(_e__�_�_�_ �_v_�_�_�_o�׻QZ_EDIT4���#TCOM_C_FG 1��'%�to�o�o 
Ua_A�RC_!"��O)T�_MN_MODE�6�Lj_SPL��o2&UAP_CP�L�o3$NOCHE�CK ?� � Rdv� ���������*�<�N�`��NO_?WAIT_L 7Jg650NT]a���Uz	���_ERR?12���ф��	���-����R�d����`O�����| ˯�
aB����o����C���������,V<� �� ?��Uϟj����قPA�RAMႳ��N�oR�=��o��� = e������ گ�ȯ��"�4��X�j�F�<�蜿��A��ҿ�"ODRDSP��c6/(OFFSET_CAR@`�o��DIS��S_A��`ARK7KiOPEN_FILE4��1�aKf�`OPTION_IO�/�!���M_PRG %��%$*����h�WmOT��E7O�����Z��  N�� �Z"�÷�"�	 �V"�Z����RG_D?SBL  ���ˊ���RIEN�TTO ZC����A �U�`IM_D���O���V�LCT �@��Gbԛa�Zd�׏_PEX�`7�*�R[AT�g d/%*�>�UP ���{������������_�$PAL��������_POS_CH�U�7����2>3�L�XL�p��$�ÿU�g�y� ��������������	 -?Qcu����Y2C��� "4FXj|� ����� //$/�6/H/Z/l/~/�Y�@��.��/�/ςP�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO �/�/LO^OpO�O�O�O �O�O�O�O __$_6_ H_Z_)O;O�_�_�_�_ �_�_�_o o2oDoVo�hozo�o�o�_<�!��o�m ���~ BPw�m�m���~�jw8��w��� ���2�T��p��w���H��t	`���̏<ޏ��:�o������ �2��pA�  I��j�`������ ���џ���@���#�)�Or�1���� 8�}��, �\����� @D�  &��?���~�?� ���!D������G��  ;�	l��	� �xJ젌����㠯 �<� ����%�	�2�H(��H�3k7HSM5G��22G���GN�3%�R��oR�d��2�Cf��a��{���������/��3��-¸��4��>����𚿬���3�A�q�½{q�!ª��ֱ� "�(«�p=�2����� ��_{  @�Њ��_�  ��Њ��2���.�	'� �� ��I� ��  �V�,�=�������˖ß���  �y��n @"��]�<߼+"������-�N�Д߇  '�Ь�w�ӰC>��C��\C߰���Ϲ��ߤ!���@%�4���/��2�~�B��B�I�;�)�j客z+���쿱����������( �� -��#�������!�]�9�|�  q�?�ffaH�Z��� ������"��8� ����>�|P$��}�(� ��P��������\�?���� x� ���<
6�b<߈;܍��<�ê<���<�^�*�gv�A)ۙ�脣��F��?fff?}�?&�� ��@�.���J<?�\��N\��)������� ����ޤy�N9 r]������ �/&/�J/5/n/��	g/�/c(G@� G@0i�G�� G}���/??<?�'?`?K?�?o?BL
i�B��A�?y?�?|� �?K�?ů�/QO�/xO��?�O�O�O�Om��bs��n�t @|�O '_�OK_6_H_�_lS��!A��RS�i�Cn_�_xj_0O�]?��o�oAo,o¹�Wi����ToC���`CH�Qo>Jd�`a�a@�Iܚ>(hA�� �ALffA�]��?�$�?����ź°u��æ�)�	ff���C�#�
ܢopg\)��3�3C�
������<��nG��B���L��B�s�����	0źH����G��!G���WIYE����C�+�½I�۪I�5�H�gMG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo�� �
��U�@�y�d��� ������я����� ?�*�c�N���r����� ���̟��)��9� _�J���n�����˯�� �گ�%��I�4�m� X���|���ǿ���ֿ ���3��W�B�Tύ� xϱϜ���������	� /��S�>�w�bߛ߆� �ߪ߼�������=��(�a�L�(q���)����Z�������a3�8�������a4Mgux�����a�VwQ��(�4p�+4�]B�B���p�����������UPbP���Q O%x�1[FjR�������  C���I 4mX�8
O������.//>/d/R/�Rj/|/�/�/�/�/�/:  2� Fs�gGT]�&6�M�eBmpX�R�P�aC��3@�_ p?�?�?�?�?�?�=�S�OO)O;OMO�c�?���@@�jJ��`�`�1�`�^
 TO�O�O �O�O�O_#_5_G_Y_�k_}_�_�_�j�A �����D��$�PARAM_ME�NU ?B���  �DEFPULS�E{	WAIT�TMOUTkR�CVo SH�ELL_WRK.�$CUR_STY�L`DlOPT�Z1ZoPTBooibC�?oR_DECSN `���l�o�o�o &OJ\n������QSSREL_ID  >��
1��uUSE_P�ROG %�Z%8�@��sCCR` ��
1�SS�_HOST7 !�Z!X����M�T _���x�������L�_TIME�b �h��PGDE�BUG�p�[�sGI�NP_FLMSK��E�T� V�G�PG�Ar� 5��?��CyHS�D�TYPE�\�0��
�3�.� @�R�{�v�����ï�� Я����*�S�N� `�r����������޿ ��+�&�8�J�s�n���ϒϻ�G�WORD� ?	�[
 	�PR2��MA9I�`�SU�a��cTEԀ���	Sd�COL��C߸��L� C�~��h�d*�TRACE�CTL 1�B���Q �� �'��0�ށ�_DT Q�B������D � �a�A�������	��
�������Y�Y�Y����Y��	0�ґ@�� �@�Ҩ��҅@������ ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9�K]�� ���������S0��� "HH�@JHU�&ЎЖОUЦЮжоU����ҎҖUҞҦҮҶUӎӖӞӦUӮӶҾ���Ҿ�����Ҫ��&�.Ҫ6����� ��hz�� ���/�/�/�/�/�/  ??$?6?H?Z?l?~? �1�ь%(O:OLO^OpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����� ����*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟڟ���� "�4�F�P�$Or����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~�f��� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo�xo�o�o�o�o�o�a��$PGTRACE�LEN  �a � ����`��f_UP _����q'p�q p�a_CFoG �u	s�a0q�Lt�ceqx>c}  �qu4r�DEFSPD e�?|�ap��`�H_CONFIG� �us ��`�`d�t��b 	�a�qP�tcq��`ۂ�`IN7pTROL �?}_q8�u��PE�u��w��qLt�qqv�`L�ID8s�?}	v�L�LB 1��y ���B�pB4Ńqv �އ؏�	�s << �a?��'��� A�o�U�w�������۟ ��ӟ��#�	�+�Y�v�񂍯����ï
���������/�u�GRP� 1ƪ��a@�j��hs�a�A�
D�� �D@� Cŀ @�٭^�t������q�p���.� ����Ⱦ´���ʻB �)�	���?�)�c���a>��>�,᷁Ϻ��ζ� =4?9X=H�9��
� ���@�+�d�O���s���o߼�����  Dz���`
��8��� H�n�Y��}����� ��������4��X�C��|���)��
V7�.10beta1�Xv A���ι��!�����?!�G�>\=y��#��{33A!���@��͵���8wA��@�/ A�s�@Ls���� ��"4FXLs�ApLry�ā���_��@l��@W�33q�`s��k��Anff�a���ھ��)7�x�� �ar� T�n�t����	�t�KNOW_M � |uGvz�SV ��z�r�&� ���>/�/G/��a��y�MM���{� ���	^r�` (l+/�/',�$�@XLs	����@���%�"�4�.N�z�MRM��|-TU�y�c?u;e�OADBANFW�D~x�STM�1 �1�y�4Garra_B�2Sem��?~s�;Co�2��O�7��3Antena�_Full @� �VODe�qH��^OpO �O�O�O�O�O�O!_ _ _W_6_H_�_l_~_�_��b�72�<�!4�_ � �<�_�_N�3 �_�_
oo�749oKo]ooo�75�o�o�o�o��76�o�o�77 2DVh�78��X���7MA�0���swwOVLD � �{�/a�2P�ARNUM  p�;]��u�SCH*� 8�
����ω�3�UPD��[�ܵ+�>wu_CMP_r -���0�'�5C�ER�_CHKQ���`�1�"e�N�`�RS>0��?G�_MO�?_���#u_RES_G
�0��{
Ϳ@�3� d�W���{�������� կ���*�����P��O��8`l��� ����`��ʿϿ��` �	���1p)�H�M� ��phχό���p��x�����V 1��5|�1�!@`y�ŒTHR_INR>0�/�Z"�5d:�MASmSG� Z[�MNF��y�MON_QUEUE ��5�6ӐV~  #tNH�U��qN�ֲ���END�����EXE������BE������OPT�IO������PROGRAM %���%��߰���TA�SK_I,�>�OCFG ά�]���^��DATAu#�����Ӑ2�%B�T� f�x���5��������������,>P�IWNFOu#� ���� ����� '9K]o��� �����/lx�� � ;���ȀK�_�����S&ECNB-�b-&q�&2�/ڝ(G��2�b+ �X,		��=�{���/��@��P4$�0��99)�N'�_EDIT ����W?i?��WERF�L�-ӱ3RGAD�J �F:A�  �5?Ӑ�5Wј6���]!֐��??�  Bz�WӐ<1Ӑn&%�%O�8�;��50!2��7�	�H��l0�,�B=P�0�@�0�M�*�@/�B *�*:�B�O�F�O2��D��A�ЎO�@O	_�,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_�_o �_o�_�_
o�o.o�o jodovo�o�o�o�o�o �o\XB<N� r����4��0� ��&���J������� ����������x� "�t�^�X�j�䟎��� ʟğ֟P���L�6�0� B���f���������(� ү$������>��� z�t��� Ϫ����� �l��h�R�L�^�DX�	���ώ0�� ���t$ :�L��o�
���ߥ��7PREF S��:�0�0
�5?IORITYX�M6}��1MPDSPV��:n" �UT��C�6�ODUCT���F:��NFOG[@_�TG�0��J:?�HI?BIT_DO�8���TOENT 1��F; (!AF�_INE*������!tcp����!ud��8�!�icm'��N?�X�Y�3�F<��1)�� �A�����0� ����������'  ]D�h�������*>��3���9n"OTf�3>�)��2�B�G/�LC���4�;LFJAB,  ���F!/�/%/7/�5�F�Z@�w/�/�/�/�3&�ENHANCE S�2FBAH+d�?�%;�������Ӓ1��1PORT_N�UM+��0����1_CARTRE�@��q�SKSTyA*��SLGS�������C�U�nothing�?�?OO�۶0TEMP �N�"O�E��0_a_seiban|߅OxߕO�O �O�O�O_�O'__K_ 6_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1U@e� v����������Q�<�u�.IVE�RSI	�L��� �disabl�e�.GSAVE ��N�	267_0H771|�h���!�/��9�:� !	^�4�ϐ����e��͟ߟ������9�D�C-Å_y� +1���������ő����Ǻ�URG�E� B��r�WF Ϡ��-��9�W�����l:WRUP_DELAY �=�n�WR_HOT �%��7��/p��R_NORMALO��V�_�����SEMI𓿹�����QSKI%Po��97��xf�=� b�a�sυ�H��ʹ��� ���������&��J� \�n�4�Fߤߒ����� �߲���� �F�X�j� 0��|�������� ���0�B�T��x�f����������ãRBT�IF�5���CVT�MOU�7�5����DCRo���� �T�C���C���C��?���>�<�h=@�jH�������=W%±�;���x$�4?s#�HG�HϘ��� <
6b<�߈;܍�>�u.�>*��<��ǪP0���2DVhz��������,GR�DIO_TYPE�  v��/ED�� T_CFG ���-�BH]�E�P)�2��+ ��B�u �/�*��/ �?�/%?=�/V?� }?�Ϟ?���?�?�?�? �?O
O@O*Gl?qO�� 8O�O�O�O�O�O�O�O �O_<_^Oc_�O�__ �_�_�_�_�_o�_&o H_Mol_o�oo�o�o �o�o�o�o�o"DoI ho*j���� ���.3�E��f�  ���x��������ҏ �*�/�N��b�P��� t�����Ο��ޟ�:��+���R'INT 2��R��!�1G;�� i�{��"���8f�0 ��ӫ��� ���M�;�q�W��� ����˿���տ�%� �I�7�m��eϣϑ� �ϵ�������!��E� 3�i�{�aߟߍ��߱߀��������A���E�FPOS1 1�~!)  x� ��n#���������� ����/��S���w�� ��6�����l����� ��=O����6�� �V�z� 9 �]����R d���#/�G/� k//h/�/</�/`/�/ �/??�/�/?g?R? �?&?�?J?�?n?�?	O �?-O�?QO�?uO�O"O 4OnO�O�O�O�O_�O ;_�O8_q__�_0_�_ T_�_�_�_�_�_7o"o [o�_oo�o>o�o�o to�o�o!�oEW�o >���^�� ���A��e� ��� $�����Z�l����� +�ƏO��s��p��� D�͟h�񟌟�'� ԟ�o�Z���.���R� ۯv�د���5�ЯY� ��}���*�<�v�׿¿ ����Ϻ�C�޿@�y�<�e�2 1�q�� -�g�����	��-��� Q���N߇�"߫�F��� j��ߎߠ߲���M�8� q���0��T���� �����7���[���� �T�������t����� !��W��{� :�^p�� A�e �$�� Z�~/�+/�� �$/�/p/�/D/�/h/ �/�/�/'?�/K?�/o? 
?�?.?@?R?�?�?�? O�?5O�?YO�?VO�O *O�ONO�OrO�O�O�O �O�OU_@_y__�_8_ �_\_�_�_�_o�_?o �_co�_o"o\o�o�o �o|o�o)�o&_ �o��B�fx ��%��I��m�� ��,���Ǐb�돆�� ��3�Ώ���,���x� ��L�՟p�������/� ʟS��w�����ϓ�3 1��H�Z��� ���6�<�Z���~�� {���O�ؿs����� � ��Ϳ߿�z�eϞ�9� ��]��ρ���߷�@� ��d��ψ�#�5�G߁� ������*���N��� K����C���g��� ������J�5�n�	� ��-���Q������� ��4��X��Q ���q��� T�x�7� [m�//>/� b/��/!/�/�/W/�/ {/?�/(?�/�/�/!? �?m?�?A?�?e?�?�? �?$O�?HO�?lOO�O +O=OOO�O�O�O_�O 2_�OV_�OS_�_'_�_ K_�_o_�_�_�_�_�_ Ro=ovoo�o5o�oYo �o�o�o�o<�o` �oY���y ��&��#�\��������?�ȏ����4 1�˯u�����?�*� c�i���"���F���� |����)�ğM���� �F�����˯f�﯊� ����I��m���� ,���P�b�t������ 3�οW��{��xϱ� L���p��ϔ�߸��� ���w�bߛ�6߿�Z� ��~�����=���a� �߅� �2�D�~����� ���'���K���H��� ���@���d������� ����G2k�* �N����1 �U�N�� �n��/�/Q/ �u//�/4/�/X/j/ |/�/??;?�/_?�/ �??�?�?T?�?x?O �?%O�?�?�?OOjO �O>O�ObO�O�O�O!_ �OE_�Oi__�_(_:_ L_�_�_�_o�_/o�_ So�_Po�o$o�oHo�o�lo�oۏ�5 1� ���o�o�olW��o �O�s���2� �V��z��'�9�s� ԏ���������@�ۏ =�v����5���Y�� }�����۟<�'�`��� �����C���ޯy�� ��&���J����	�C� ����ȿc�쿇�ϫ� �F��j�ώ�)ϲ� M�_�qϫ����0��� T���x��u߮�I��� m��ߑ�������� t�_��3��W���{� �����:���^���� �/�A�{����� �� $��H��E~� =�a����� D/h�'�K ���
/�./�R/ ��/K/�/�/�/k/ �/�/?�/?N?�/r? ?�?1?�?U?g?y?�? O�?8O�?\O�?�OO }O�OQO�OuO�O�O"_<t6 1�%�O �O_�_�_�_�O�_|_ o�_o;o�__o�_�o o�oBoTofo�o�o %�oI�omj� >�b����� ��i�T���(���L� Տp�ҏ���/�ʏS� �w��$�6�p�џ�� �������=�؟:�s� ���2���V�߯z��� ��د9�$�]������ ��@���ۿv�����#� ��G�����@ϡό� ��`��τ�ߨ�
�C� ��g�ߋ�&߯�J�\� nߨ�	���-���Q��� u��r��F���j��� ����������q�\� ��0���T���x��� ��7��[��, >x����!� E�B{�:� ^�����A/,/ e/ /�/$/�/H/�/�/ ~/?�/+?�/O?5_GT7 1�R_�/?H? �?�?�?�/O�?2O�? /OhOO�O'O�OKO�O oO�O�O�O.__R_�O v__�_5_�_�_k_�_ �_o�_<o�_�_�_5o �o�o�oUo�oyo�o �o8�o\�o�� ?Qc���"�� F��j��g���;�ď _�菃������ˏ� f�Q���%���I�ҟm� ϟ���,�ǟP��t� �!�3�m�ί��򯍯 ���:�կ7�p���� /���S�ܿw�����տ 6�!�Z���~�Ϣ�=� ����s��ϗ� ߻�D� �����=ߞ߉���]� �߁�
���@���d� �߈�#��G�Y�k�� ���*���N���r�� o���C���g����� ������nY�- �Q�u��4��X�|b?t48 1�?);u�� /;/�_/�\/�/ 0/�/T/�/x/?�/�/ �/�/[?F???�?>? �?b?�?�?�?!O�?EO �?iOOO(ObO�O�O �O�O_�O/_�O,_e_  _�_$_�_H_�_l_~_ �_�_+ooOo�_soo �o2o�o�oho�o�o �o9�o�o�o2�~ �R�v���5� �Y��}����<�N� `���������C�ޏ g��d���8���\�� ��	�����ȟ�c�N� ��"���F�ϯj�̯� ��)�įM��q��� 0�j�˿��ￊ�Ϯ� 7�ҿ4�m�ϑ�,ϵ� P���tφϘ���3�� W���{�ߟ�:ߜ��� p��ߔ���A�����  �:����Z���~� ����=���a����� �����MASKW 1����������XNO  ����� MOTE � �R_CFG� �Y����P?L_RANGUP�����OWER ���� �A���*SYSTEM�*P�V9.304�4 �1/9/2�020 A ��� ���REST�ART_T  � , $FLA�G� $DSB_�SIGNAL� �$UP_CND�4� �RS232�r � $�COMMENT �$DEVI�CEUSE4PE�EC$PARIT�Y4OPBITS�4FLOWCON�TRO3TIME�OUe6CU�M�4AUXT��5INTERFACs�TATU� �KCH t $OLD_y�C_SW 'F�REEFROMS�IZ �ARGE�T_DIR �	$UPDT_M�AP"� TSK_wENB"EXP:*z#!jFAUL �EV!�RV_D�ATA�  �$n E�   �	$VALU�!� 	j&GRP_ �  {!A�  2 �S�CR	� ��$ITP_�" �$NUM� OU�P� �#TOT_A�X��#DSP�&J�OGLI�FIN�E_PCd�ONmD�%$UM�=K5 _MIR1!4�PP TN?8APL"G0_EXb0<$�!�� 814�!PGw6BgRKH�;&NC� �IS �  �2T�YP� �2�"P+ Dxs�#;0BSOC�&�R N�5DUMMY�164�"SV_C�ODE_OP�S�FSPD_OVR5D�2^LDB3�ORGTP; LEbFF�0<G� OV5;SFTJRUNWC!�SFpF5%3UFR�A�JTO�LCH�DLY7RECO1VD'� WS* �0��E0RO��10_~p@   @��}S NVERT"�OFS�@C� "F�WD8A�D4A�1EN�ABZ6�0TR3�$1_`1FDO[6MOB_CM�!FPB� BL_M��!2hRnQ2xCV�"' } �#2PBGiW|8AMz3\P0��U�B�__M�P��M� �1�AT$CA�� �PD�2�PHB�K+!:&aIO�4 �eIDX+bPPAj?a$iOd7e�U7a��CDVC_DBG "�a;!&�`�B5�e�1�j�S�e3�f�@ATIO� ���AaU�c� �S�AB
0Y.#0�D��X!�� _�:&SUBC�PU%0SIN_RS�T, 1N|�S�T�!�1$HW_C�1�"]q.`�v�Q$�AT! � �$UN�IT�4�p�pAT�TRI= �r0CY{CL3NECA�b�L3FLTR_2_�FI9a7�c,!L�P;CHK_�S�CT>3F_�wF_�|8��zFS+�R�rCHAGp�y��R�x�RSD�@'�1E#�&7`_T�XPRO��`@S�EMPER�_0�3Tf�]p� xf��P�DIAG;%?RAILAC�c4r�M� LO�0�A�65&�"PS�"�2 -`�e��SPR�`S.  ��W�Ctaf	�CF�UNC�2�RINS_T.!(�w�L�� S_� �0�Pp�� 	d��WARL0~bCBLCUR���єAʛ�q͘ƘDA`�0���ѓʕLD  @,a3��!��8�3��TID�S��!� $?CE_RIA !5+AFDpPC~��@��T2 �C9#�b{Q�OI�pCVDF_LaE��#0(!�LM�S�FA�@HRDYO,L1	PRG8�H��>1�(�ҥMULSE� =#Sw3��$J�JJ6BKGFKFAN?_ALMLV3R��WRNY�HARDH�0+&_P "��2Q�Ȏ�!�5_�@:&AU��Rk��TO_SBRvb��� ƺ�pvc|�޳MPINF�@��q�)���REG�'d~0V) 0R�C�1DgAL_ \2FL�u�2$MԐ(�#S�d�P� `�g�CMt`3NF�qsONIP�q�E�IPP 99a$Y��!� �"�!� �o3EGP��#@F��AR� �c�52������|5AXE�'R�OB�*RED�&W�R�@�1_=��3SYР0ѥ0_�Si�WR1I�@�ƅpST�# ��0*@� �q	���3���� B� �A��3�D.�POTO�� �@ARY�#��!��d�!�1FI�0�$LwINK��GTH�MB T_���A��96�"/�XYZ+"9�7G�OFF�@��.�"���B� l�`���A3$ ��FI�p����4�4l��$_Jd�"(B�,a������8�"q������Ck6DUR��9.4�TURT�XZ�N�����Xx��P��FL�/�@s��l�P��3y0�"Q 1� %K
0M:$�53]q7�pSuD�Sw#ORQɆ@�!�����Q7��0O[ЁND�=#�!#�1OVE8��M��� R��R��Q!P.!P! OAN}q	�R ����990� �brJ�9V����v�!E)R1��	8�E�@n $D�A��p�嘕`Ă���v�AX�C �"��`�q�s� ��0~3�~F�~@e�~�~E�~1�� ~Ҡ{Ҡ�Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�Ҡ��Ҡ�!)DEBU}s$x���삼!R*�AB�a8A29V`|r 
�"�c ���%�Q7�7�17 3�7F�7e�7�7�E�������LA�B����yp�cGR�O�p��}��PB_ ҁ ��̓��ð�6�1p���5���6AND���8p�a3���-G  �Q����AH�PH�p2��NTd��Cs@VEL�؁�}A��F�SE�RVEs@�� $�����A!�!�@PAOR}�KP�иA�Bl���	��$�BTRQ�
�CH��@
�G��2	�Eb��?_  lb��QN�ERR��RI�P8�@�FQTOQ�� AL�}��YVĀG�E�%�\ ���ARE>�  ,�A�E�P
�RA�Q O2 d�R7c�Un�@ ��$F �ׂ��m �COC|��P  8[�COUNT�ђSF�ZN_CFG�A# 4�p%��rT\zs �a�#`pJp�qY�&c��/ �� MGp+�����`�OGp�eFAq����cX8еk�i�oQ��'ѴDp8�P�z��@HELA�-b� 5��B_wBAS\RSR$Ɗ`�2�S��L�!p1T�W!p2Dz3Dz4DzU5Dz6Dz7Dz8�WqROO���P�1�3NL�� �AB�C
�n"pACK�&IN�P	T+�W�U��	�k��y�_PU8�~�|�OU�CP��%�s�Vl����YTPFWD_KcARKQ-�:PRE�D��P����QUE�$�Ā9 )���~���I U��#s/���@�/�SEM1ǆ1�An�aSTY�tSO����DI�q��Qc��X_TM9�MANsRQ �/�END���$KEYSWI�TCH2�G����H}E)�BEATMz�PE��LEJR���0Jx�UF�F��G�S��DO_HOM��Olz��pEFPR��PSbJі��uC��O��<7P�QOV_M��}�c�IOCM���1��� uHK�� �D,�&�a`U2R��M���a�r +�FORC�*�WAR��OM>��  @�$��*��U��P�1��g����3��4�1�B�PO�W�Lz��R%�UN�LO�0T�ED���  �SNP���S.b 0N�A�DDa`z�$SI=Z*�$VA�0�U�MULTIP�r����Az� � $��ƒ����SQc�1CFPv�FRIFr�PSw���ʔ�f�NF#�ODBU x�R@w������F��:��IAh�����������S"p�� � � �cRTE���SKGL.�T�x�&C`�Gõ3a�/�STMTd��`�P����BW9 �0�SHOWh�qBANt�TPo���E�����PV_�Gsb �$PC��0�PoFBv�P��SP��A�p�ş@�VD��rb�; �+QA002D.� ��6ק�6ױ�6׻�6�U54�64�74�84�94�A4�B4و�6��17�}�6�F4� �؀@�����Z����t�1���1��1��1��1���1��1��1��1���1��23�2@�2�M�2Z�2g�2t�2���2��2��2��2���2��2��2��2
��2��33����M�U3Z�3g�3t�3��U3��3��3��3��U3��3��3��3��U3��43�4@�4M�U4Z�4g�4t�4��U4��4��4��4��U4��4��4��4��U4��53�5@�5M�U5Z�5g�5t�5��U5��5��5��5��U5��5��5��5��U5��63�6@�6M�U6Z�6g�6t�6��U6��6��6��6��U6��6��6��6��U6��73�7@�7M�U7Z�7g�7t�7��U7��7��7��7��U7��7��7��7�٭7��AT��Pv�U�B �@�09r�
B�V���A x� �0R���  ��BM�@RP�`�4Q_�PR�@[U�AR��D�SMC��E2F_qU��=A�YSL�P>�@ �  �ֲ >g�������iD��VALU>e�pL�Az�HFZAID_L����EHI�JIh�$F�ILE_ ��D�d�$Ǔ�PXCSA�Q� h�0!PE_B�LCKz�.RI�7XD_CPUGY!�GY��Ic�O
T�`Y.��R�  � PaW`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q��TJ��U�Q�T�Q�UH���T`�T ��T2L�_LIz��  �pG_O�T�P_EDI�U�,/`�`7c �?bة�pBQh��� ��TBC2 �! ��%�>��P��a�7aFqTτ�d݃TDC�PA�N`�`M�0�f�a&�gTH��U��d�3��gR�q�9�ERVAEЃt݃t	��a��p�` "X ;-$EqLENЃRt݃Ep�pRAv��Y@�W_AtS1Eq�D2&�wMO?Q�S���pI�.B�A�y�4Ep�{�DE�u��LACE� �CCC�.B��_�MA��v��w�T#CV�:��wT,�;� Z�P���s�~��sёJ耭0��M����JH���uā�uQq�2ѐ���݁�s�JK��VK�������	���J����JJv�JJ�AAL�@<��<�6��:�5�cm�N1a�m�,��D�L�p_\�Ű	 v�aCF
�# `�0GROU�@J�Բ���N�`C^�ȐREQ�UIRrÀEBU�u�Aq��$T�p2�"��Bp薋a	��d$� \?@qhAPPR���CLB
$H`NN;�CLO}`K�S�e�`��u
�aI�% �3�M�`�l��_MG񱥠C �"P�����&���BRK��N�OLD����RTM!O6a�ޭ��J6`�P>��p��p��pZ�(�pc��p6+�7+�<���d�e&� ��lr��������PATH��������qxȪ����%0A��SCaAub��<���INDr�UC�p�q�C�U%M�Y�psP�����A q/ʤ�/�E�/�P�AYLOA�J2=L�0R_AN�apÁL�Pz�v�jɆ���R_F2LSHRt��LO{�R������>�ACRL_�qŐ����b��H�@B�$H��"�FLEX�>��aJ�f' P (��o�o+R?�Du( :Qcv�p ����f��po��|F1���-������]�E��*� <�N�`�r�����4�Q� ������A�c���ɏۏ$���T��2�X:A�� �������� )�;�?�H�6�Z�c�u�臟����J��) ���`��˟ݟ�`�0ATF�𑢀EL��(aj��J�(��JE۠gCTR��A�TN�1��HAND_V�BB>ѯ@�* M$��F2���d�C�SW����+� $$M�����0ˡ�@ڡ������A�@ g����A)��A���@
˪A٫A� ��`P�˪D٫D�PȰG�P�)STͧ�!ک�!N�DY�P9���� #%��Fp���Ѫ���i� ���������P3�<� E�N�W�`�i�r�����, ��ԓ� �n�5m��1ASYM$ص.@�ض+A������_`��	����D�&�8�J�\�n�J�u�&��ʧC�I��S�_�VIo�Hm��@V_UNVb�@
S+��J�"RP5"R��&T�� 3TWV�͢���&���$�U��/�7� �`�`3HR`ta-��QLQ�1�DI��O�T8�R�P��. ; *"IAA*���$aG�2C�2cJ�$?pI��P �/ � �MEB�� Mb�R4AT�PPT�@� ��ua����AP�l@zh�a�iT�@��� $DUM�MY1E�$PS�_D�RF��P$��f3�FLA��Y�P���b}c$GLB_T��Uuu`1�py���EQa0 X(����ST����S�BR�PM21_V���T$SV_ERb��O_@KscsCLp�KrA��O'b�PGLv�@EW��1 4���a$Y,Z,W�s怯��AN`¥���qU�u2 ��N��p�@$GIU{}$�q 1u8�q�p��3 L���v�^B}$F^BE�vNWEAR��NK�F8����TANCK⥑JsOG��� 4� $JOINT����� �sMSET.��5  �wE�H�� S��� ��6��  MU��?����LOCK_F�O����PBGLV�HGL�TEST�_XM>���EMP�t����r̀$1U�Гr��22���sB,�3���Ҁ,�1Mq�CE���sM� $K�AR��M�STPD�RA�pj�a�VECX��{�e�IU,�41�{HEԀTOOL�ڠ�V�RE��IS�3����6N�A�AC)H���5��O�}cj�d3���pSI.��  @$RAI�L_BOXE���ppROBO��?�~pqHOWWAR*�x��`�ROLM�b B���S��
�5����O_F� !ppHOTML5�Q��h���SGU�CH��]7m�	�R��O�ҡ8���v�z���_;OU��9 tpp(��14A�̀��PO�֡%PIP��N ��
�ڑS�,�����?CORDEDҀްL̠5�XT��q)Hb�P� O4` : 7D pOBP!" Ҁ{�j��cpj�^@$wSYSj�ADR#��Pu`TCH� 7; ,��EN�RZ�Aف_�t״�c��PVWVAPa<� � p��r�UP�REV_RT]1�$EDIT�VSHWR�7v;���J�q�@D_`#R�~+$HEADoAh�Pl�A$�KE�q��`CPSPD��JKMP��L�U�R��Fd=r�O�϶I�5S#CiNE��$�_TICK�AM���q��HN-q�> @t������_�GP��[�STYѲ�LOq���Ҫ�?�
�Gݵ%�$���t=7pS !$Q��da�e!`�f9P�0�SQUd� �<�b�ATERCy`,zuS�@ �p�Cp����d�%Oz`mcO�IZ�d�q�e�aPRM��a8�����PUQH�_DO�=�ְXS��K�VA�XIg�f�1�UR � ��$#�Е��� Y_����ET��Pۂ����5f�F�7g�A��!�1�d9�2�;�SR|Al�о���#�� 5��#��#�)#�) i�>'i�N'i�^&{��� �){����2��C�����C��WOiO{O�D�QS�SCp B h�ppDS(�k��`SPL`�ATL �I����¼bADDRE�S��B'�SHIF���"�_2CH#r��I&p��TU&p�I� C͢CU�STO��IaV��I�bDȲ,��0
��
��V�X�R`E \�����f�7���tC�#	���F���irt�TXSCR�EEl�F�P��T�INA�s�p��t̈`��Q_��0G T��fp,⧱eqBp&�uᦲu�$#�RRO�'0R���}�!��#��;UE��H ��0��r�`S�q��RSMЂk�UV����V~!�PS_�s�&C�!�)�'C��Cǂz"� 2-G�UE�4Ibvr\�&8�GMTjPLDQ���Rp����B�BL_�W�`aJS �f�>2O�qJ2�LE�U3"�T4RwIGH^3BRDxt��CKGR�`�5T�W��7�1WIDTH��H������a��7�UIu�EY��QaK d�p��A�J�
�=4�BACKH��b4�5|qX`FOD�G�LABS�?(X`I<�˂$UR(�9@����0^`H4! L 8�QR�_k��\B_`R�p͂����a^�RIAO�aM��w�0Uj0�CRۂM�L�UM�C��� ERVH��p�0P<��4NV`��GE=B#���]�&t�LP�E��E��Z)Wj'Xz'XԐ&YU5$[6$[7$[8	R����3�<���fԑ�ŁS��M�1US=R�tO <��^`1U�r�rFO
�rPRI��m����P�TRIP�m�oUNDO��P�p���`m�4�l��8#���� QWB�P.7�G s�Tf�HL�RbOS�agfR��:">c��.qR��s�~��b*�c�#�UQ.qS��o�o�#R)�>cOF�F���pT� �cOp 1Rppt/t-SppGU��P.q��pJsETw�1SUB*�� f�E_EXE���V��>cWO>� �U�`^g��WA�'��P�q!@� V�_DB�s�p��PT��`
�V�Q�r��O9R��uRAU��t�T�ͷ�q_���Ws |%�͸OWNA`>޴$SRCE � ��D��\��MPFqIA�p��ESPD������C���Gƒ 8)�5��!X `�`�rr޴��COP�a$��C`_w������rCT�3�q����q�����@� �Y"SHADO�W�ઓ@�_UNS�CA��@��4M�DGyDߑ��EGAC��,S�PPG�Z (0NO�@�D<�kPE�B��VW�� �G���![ � ���VEE#�aڒANG�$��c薴cڒLIM_X�c��c � ����#��`� ���bVF� �s�VSCCjв�\ՒC{ЃRAlצ���RpNKFA��%�E���Z`G� ^0[��C`DEĒ��� STEQ1���@�ꁻ@ I��`+0����`����P_A6�r���K�|���!]� 1�������\��сCP9C�@]�DRIܐ\�B͑V#Ѐ���D�T?MY_UBY�T��@�c��F!���Y�브����P_V�y��L�N�BMQ1$��DEY��EX�e���MU��X�M� U1S�!���P_R��b��P� ߖG��PACIr�ʐf�ᔟ��c���c���#�EqB��a�WrB����^ ܀GΐP����`C�R~``�_�0�@3!��1zr	�e�R�S�W��p�Yp��S�6�OD�Q�1A� X�#�E��UE��Yp)�D�HKJ�`�@p���8U� �EAN�ٖp��pXՆ`C�MRCV��!a ��@O��M
�pC�	��s����REF*7
������ ��/��P��@���@��b��֗�_Y��ژ��� ���Q$3����Ӷ�C��$b ����%����Q��$GRO�U� �c�����ʠ]��I2^0��U` 0_�I,�o � +ULա`��C&�rA3aB�?�NT���􀲂���A���Q��K�L ����õ��A���Q���T a$c t�`MD�p8�HU����SA�CMPE FP  _�Rr��p@����XS	��V�GF/�b#d, �&�@M�P^0۰UF�_C !���z �RO h0"+���@���0C��UREB���RI��
IN�p������d��d��ca�IN"E�H�y��0V�a-�걗�3�W����`���C��i�LO��}�z�@0�!�QNSI��݁���c$&�c$&^.�X_PE-YW+'Z_M�ڒW�Iӑ$�" �+R�'rR;SLre �/�IM
`�RE�C7�Gd�۰�̵ҭ�q��� �u��Ȑ���`���S_P�VnP ���IA�vf �~pHkDR�p�pJO�P���$Z_U�P��a_LOW��5�1J�dA��LINubEP?�tc_i�1H�1���@�G1@m�0|W�xg 5X�PATHP X�CACH$�]E��PyI�A��{�C�ID3�FA�ETD�H��$HO�pO�b@�{��d6�F�����p�PgAGE�䁀VP��<��(R_SIZ��2T�Z3�-X�0U�q�M�PRZ��IMG����AD�Y�MRE��R7WGP��8�p���ASYNBUF�VRTD�U�T7Q>�LE_2D-��U���`CҡU1��Q�u��UECCU��V�EM��]EDb�GVIRC�Q�U�S�B�Q��LA��p�NFOU�N_�DIAG�YR�E�XYZ�cE�W@Ѵh8�dpqa`T��2�IM�a�V|be��E_GRABB��Y�.a�LERj�C4���1FC-A�6504x��D7u����V���h��}`�CKLAS_@pl�BA��N@i  G��T��� @ݲմ$8BAƠwj �!q�eb��uTYSp�H�����2��I�t:b�f��B�)�EVE����PK����fx��GI�pN�O��2� \r_HO|����k � �� �
8�Pi�S�0ޗ���RO�ACCEiL?0=���VR_�U7@�`��2�p��A�R��PA��̎K�D���REM_But �D�rJMX �l|�t�$SSC�U�k@C�0G�QN@m I� �S�P�NS���VLEX�vn{ T�ENAB x2�W@��FLDRߨFI�P�t�ߨ(Ğӽ�0�VP2HFoO� ��V
>Q MV_PI��@8T@󐉰�F@�Z�+�#��8��8#��GAB���LsOO��JCBx���w"SCON(P�P�LANۀ�Dp�3F �d�v�9PէM��Q ;����SM0E�ɥ� 8ɥWb72$`<�8T���,`RKh"ǁV�ANC���R_Ou N@p (�-#<#pc��c2�w�9A/�N@q 4�������`	�^�� w�N@r� hn���1^�&OFF`|�p�`��`��DEA�
�P,`SuK�DMP6VIE���2q q �a���rs < {���4����r{7��D���^L�CUST�U���t $G�TIT>1$PR\���OPTap ��VS)F�йsu�p�0`rt&�@ASMOw�vI�|�ĄJ����%�eQ_WB��wI����� @O3�@�XVMRxxmr��T��C�ZABC��y op����)��
t�ZD$�CSCH��z Lu����`��2�%PC ��7PG�N ��<��A��_F�UNH��@��ZI�Pw{I��LV�,SL��~���Z/MPCF��|��E�����X�DMY_L�NH�=�D�� ��} $�A� ]�CMCM� C,SC�&!��P�� '$J���DQ��@�����������_�Q�,2����UX�a\�UXEUL��a�������(�:�(�J���F�TFL��w��Z�~Zp+�6����Y@Dp � 8 $R�PU<��> EIGH����#?(�iֱ�b���et� �a����У$B�0�0@�	�_�SHIFD3-�RV2V`F�@��	$5��C�0��&!�������b
�sx�uD�T�R��V̱_��SsPH���!� ,���������4A�R�YP��%������%���"�%! U �H�(UN0 ���"�2������K��q0GSP1Dak����P ��O����0���ֱ�"!NGwVER`q i�w+I_AI�RPURGE  =i  i/��F`E�Tb� �+ � � h2ISOLWC  �,�"�!D!�%��P+�_/�*OB��Dm�?�@�!H771  34n?�?@�9� `�E/#�)x� �S232�� 1�i� LT�Ek@ PENDA`�341 1D3<�*? Ma�intenanc�e Cons B��? F"O,DNo UseMJOOnO��O�O�O�O2�2NPQO;� 19%�1;CH=� �-Q�		9Q_!U�D1:___RSM�AVAIL/�/%��A!SR  ��+��H�_�P1�TVAL.&���P(.r�YVL�}� 2i��� D��P 	�/_oUQNo�orc i�o�g�o�o�o�o�o *,>tb� �������� :�(�^�L���p����� ��܏ʏ ��$��H� 6�X�~�l�����Ɵ�� �؟�����D�2�h� V���z��������ԯ 
���.��R�@�b�d� v�����п��������(�N�<�r�i�$�SAF_DO_PULS. jQp��F��CA� �/%�&�0SCR �`X�_�0�0�
	14�1IAIE���b vo$�6�H�Z�l� ~�ߢߴ���������V�HS��2%�D��d1�(�8�rb��� @�"k�}��T�h� J`����_ @��T�7 �����#�0�T D��0�Y�k�}� �������������� 1CUgy�O�Ef�����  �5;��o�� 1p�U�
�t��Di��������
  � ��*������gy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�?��?�?OO%O7O<A� ��`OrO�O�O�O�O�O �O�O?O�_._@_R_ d_v_�_�_�_�_�Q _�R0MJTo!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏJO ��'�9�K�]�o��� ����_ɟ۟���� #�5�G�Y��_�U�_�� ������ϯ���� )�;�M�_�m������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T�f�;�?�q߮��� ��������,�>�P� b�t�������������������Y��	12�3456781�h!B!����F������� ����������  ��;M_q��� ����%7 I[l*���� ���//1/C/U/ g/y/�/�/�/n��/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O �/)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_O_�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�op_�o �o�o/ASe w������� ��o+�=�O�a�s��� ������͏ߏ��� '�9�K�]�������� ��ɟ۟����#�5� G�Y�k�}���������s�կ�w����0�L�CH  B}pw�   �=��2�� }� =�
���  	�o�ί��ǿHٿ���r������ @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖ�%Ϻ����� ����&�8�J�\�n� ��������������"�Q�*�����;��<M���D���  �]�w�*�Z�|����t  d�����*�`*��$S�CR_GRP 1�*P3� �� �*�� 6�	 _�
 ��<�+*�'U8C|@��y�yD� W�!�y��	M-10i�A/7L 1234567890���� 8��MT� � �
�	L��Y	Č� N
����Y���y�
M_	P������ ,��H�
 ���1/@@A/g/y/H�ߙ!T/��/P/�/3��+���/B�S��,?*2C4&9Ad�R?  @s�j5N?�7?��7&2R��?�}:&F@ F�`�2�?�/�?�?OO -OSO>OwObO�O=j1��2�O�O�O�O�DB� �O�O;_&___J_�_n_ �_�_�_�_�_o�_%o��5j�eSgxo6����uo�o�b�1�B�|�3�oh0�4j9j9B� w�$Y̯@�HtA�Nhcu�/�%$pp�drsq ����z�q�x� �� (&�*�2�D��V�oz�e�������ECLVL  ��g��iqpQ@���L_DEFAUL�T ���s�փHOTS�TR�qq��MI�POWERF��xH���WFDO�� �RVEN�T 1ɁɁ�� L!DUM_�EIP�����j!AF_INE�<����!FT}�֞�����!-/� ���F�!RPC�_MAING�)��85���Y�VISb�t�y���ޯ!TPѠ�PUկ��dͯ*�!�
PMON_PR'OXY+���e�v���D���fe�¿!RDM_SRVÿr��g���!R,d*ϑ�h��Z�!
[��M����iIϦ�!?RLSYNC�����8����!RO�S|���4��>�!�
CE�MTCO�M?ߓ�k-ߊ�!	�S�CONS�ߒ�l�y���!S�WAS�RCݿ��m��"�!�S�USB#n|�n�!STMC��o]�����ѳ�����,���P�V�I�CE_KL ?%�d� (%SVCPRG1S������2�������o����4�������5��6;@��7ch��$���9����%� �������0�� ��X�����-� ��U���}���  /���H/���p/�� �/��F�/��n�/ ��?��8?��� `?��/�?��6/�?�� ^/�?��/X�j��q� ��#OhO��lO�O{O�O �O�O�O�O�O _2__ V_A_z_e_�_�_�_�_ �_�_�_oo@o+odo Oo�o�o�o�o�o�o�o �o*<`K� o������� &��J�5�n�Y���}�एȏ���^�_DE�V d���MC:�4��~�GRP 2d��
@�bx 	_� 
 ,V�
@�s�Z������� �����ߟ��@�'� 9�v�]�������Я��P��۫Y��
@� ܯ�P�7�t���m�����οӱ����	�� -��Q�c�Jχ�nϫ� ��X�!��ϡ��ߡ� K�!�^�p�Wߔ�{߸� �߱��������6�H�/�l���]�
y��^� ���������%��I� 0�Y��f�������� ��������3��T7]�e�����) ��
�.@�d K�o���Q����!/G/��� R/�/�/�/�/�/"�/ �/??C?*?<?y?`? �?��?�?�?�?�?�? -OOQO8OaO�OnO�O �O�O�O�O_�O)_;_ "___�?�_�_L_�_�_ �_�_�_o�_7oo0o moTo�oxo�o�o�o�o �o!x_E�oU{ b������� �/��S�:�w�^�p�𭏔�я�d �X��ZI6 r �	 @Z���0�+A�����dBjBA�=��������B���AZ.��AĊ�+ߓA.�Q�B�����5\��i�6�A�u��?'���%�����%PEGA_�BARRA_ES�TEIRA�����X�T���?=���=X��7
��?�>�A�����������&���������AxP���f��U�'A��j��´��B�:�<��3����jB]+��T��C%�T���d�ʐ����>�pc?��7��ԳT@6���A�_��0n�����·��Ak��۸I��K9FA�G�����B!v,��-��C3������pBM�@>�#�b�(�Y��������HX�?L!����Q�B����AJ��Xk��@fD3��O��A����ݒ��Yw����.B�B�;���CH�z�B�?���6����-Ϙ�����n���=]���V�@�?,߱��Ö� �����eAk�������OYߠA�ㇾ��A�B�J�;%��C$4�aƿBXZ9���
����ߘ�Ţ�� ����(��^_��-\¯ԡ��گ���+���������h���ߔ�ᢧ��*���6�>�ԯb����zװ
��BM��s��x�����U<�߯7@6|=����$�6�j�� N�@���b�G���L�}�������x7��~K@����V�+A>r�rF���������Y@�+�@�<B��|ߞA�F�����B)��,o��?ɇ��~0��0~6�Z� �Q�杚��������Aߍ��]ܖA����������2[�����>�ȥ�A��=�³�N�B �$�w�?�dj��to�7\�
�.��%��Z�����A�����*��@Ve�B� ������YN��#�BD��	���9�A���gB�#
q�3��C�4#��,?[B�VM���C�OLOCA_PR�ENS���X�\{B*3Vhz �������/
% ���/�/??B?0? R?x?�?f?�?�? �?�?OO(O~?�?uO �?NO�O�O�O�O�O�O _VO;_zO_n_ _~_ �_�_�_�_�_._oR_ �_Fo4ojoXozo�o�o �oo�o*o�oB 0fTv��o� �����>�,�b� �����R�t�N���� ����:�|�a���*� �����������ܟ� T�9�x��l�Z���~� �������,��P�گ D�2�h�V���z���� ��(�¿�
�@�.� d�Rψ�ʿ���x��� t�����<�*�`ߢ� ����Pߺߨ������� ��8�z�_��(�� �����������R� 7�v� �j�X���|��� ������������� 0fT�x���� ��,b P����v�� /�//(/^/��/ �N/�/�/�/�/ ?�/ ?f/�/]?�/6?�?~? �?�?�?�?�?>?#Ob? �?VO�?fO�OzO�O�O �OO�O:O�O.__R_ @_b_�_v_�_�O�__ �_o�_*ooNo<o^o �o�_�o�_to�o�o �o&J�oq�: \6�����"� dI���|�j����� ��֏ď��<�!�`�� T�B�x�f�������ҟ ���8�,��P�>� t�b���ڟ �ѯ��� ��(��L�:�p��� ��֯`�ʿ\�ڿ �� $��Hϊ�oϮ�8Ϣ� ���ϴ������� �b� G߆��z�hߞߌ��� ������:��^���R� @�v�d���� ��� �������N�<�r� `�������������  J8n��� ��^������ F�m�6�� �����NtE/ �/x/f/�/�/�/�/ �/&/?J/�/>?�/N? t?b?�?�?�?�/�?"? �?OO:O(OJOpO^O �O�?�O�?�O�O�O_  _6_$_F_l_�O�_�O \_�_�_�_�_o�_2o t_Yoko"oDoo�o�o �o�o�o
Lo1po�o dRtv���� $	�H�<�*�`�N� p�r������� ��� ��8�&�\�J�l� 菹������ڟ��� 4�"�X������H��� D�¯�֯���0�r� W��� ���x������� �ҿ�J�/�n���b� Pφ�tϪϘϺ���"� �F���:�(�^�L߂� pߦ������ߖ߸ߒ�  �6�$�Z�H�~��ߥ� ��n�����������2�  �V���}���F����� ����������.p�U ���v���� �6\-l`N �r����2 �&/�6/\/J/�/n/ �/��/
/�/�/�/"? ?2?X?F?|?�/�?�/ l?�?�?�?�?OO.O TO�?{O�?DO�O�O�O �O�O�O_\OA_S_
_ ,__t_�_�_�_�_�_ 4_oX_�_Lo:o\o^o po�o�o�oo�o0o�o $H6XZl� �o���� �� D�2�T������z� ԏ����
�@��� g���0���,���П�� ����Z�?�~��r� `�������̯���2� �V��J�8�n�\��� ����ȿ
��.���"� �F�4�j�Xώ�п�� ��~Ϡ�z�����B� 0�fߨύ���V��߮� ��������>��e� ��.��������� ���X�=�|��p�^� �����������D� T���H6lZ�~ ������ D2hV���� |��
/�/@/./ d/��/�T/�/�/�/ �/?�/?<?~/c?�/ ,?�?�?�?�?�?�?O D?)O;O�?O�?\O�O �O�O�O�OO_@O�O 4_"_D_F_X_�_|_�_ �O�__�_o�_0oo @oBoTo�o�_�o�_zo �o�o�o,<�o �o��ob���� ��(�jO����� �������܏ʏ �B� '�f���Z�H�~�l��� ����؟���>�ȟ2�  �V�D�z�h������ ׯ���
���.��R��@�v�������n�  ��$SERV_MAIL  �����ʴOUT�PUTո��@ʴRV 2�j�  � (r����
��=�ʴ�SAVE���TO�P10 2�� d 6 r Ʊ���϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>��P�b�t�����n�YP�Y��FZN_CF�G f���=��J���GRP� 2��g� ,�B   A �D�;� B � � B4=�RB{21I�HELL��f�e�)�*�=������%RSR ������& J5G�k�������.�  ��/>/P/"\/ �X/z"{ S�U'&"2�dh,�g-�"EHK 1S �/�/�/�/ #?L?G?Y?k?�?�?�? �?�?�?�?�?$OO1O�CO?OMM �S�ODFTOV_�ENBմ�e��"O�W_REG_UI��O�IMIOFW�DL~@�N�BWAIT�B�)��V���F�YTIMn�E��G_VA԰|_�A_UNIT�C�~Ve�LC�@TRY��Ge�ʰMON�_ALIAS ?5e�I%�he��o o&o8oFj�_io{o�o �oJo�o�o�o�o�o /ASew"�� ������+�=� �N�s�������T�͏ ߏ�����9�K�]� o���,�����ɟ۟� ���#�5�G��k�}� ������^�ׯ���� �ʯC�U�g�y���6� ����ӿ忐����-� ?�Q���uχϙϫϽ� h�������)���M� _�q߃ߕ�@߹����� �ߚ��%�7�I�[�� ������r����� �!�3���W�i�{��� 8������������� /ASe��� ��|�+= �as��B�� ��/�'/9/K/]/ o//�/�/�/�/�/�/ �/?#?5?�/F?k?}? �?�?L?�?�?�?�?O �?1OCOUOgOyO$O�O �O�O�O�O�O	__-_ ?_�Oc_u_�_�_�_V_��_�_�_ooc�$�SMON_DEF�PROG &����Aa� &*SYST�EM*obg �$JO0dRECA�LL ?}Ai �( �}xyz�rate 61=�>10.109.�3.46:138�64 .*�o4 �a 4 �a�o�o�ov	v}
�e11 �o �o�o]o�u�o. @R����(� �a�s����*�<�N��ߏ���7cop�y frs:or�derfil.d�at virt:�\tmpback�\��ӏd�v���}.��mdb:*.*�2���L�ݟ���2�x�:\��'���4A Пa�s����3�a%�7�ʏۯ���� $���H�	�k�}����� =�ƟX����� ��� D�ֿg�yό���/�¯ T����ϊ��.����� c�u߇ߚ�5߾�P��� ���ϫϸ�N�_�q� ���'�9�������� �&߯�J�[�m���� ��?��߉������"� ��F���i{���1@��V����� ����]o�����4748��L��/��tpdisc 0�8 ��\/�n/�/tpconn 0'�4/F/X/��/�/>��:pi�ckup_bar�ra_estei�ra.tp��em�p���[?m??<|?/0torno9?��/�?�?�?5�6lace�?�?��?dO�vO�O};�5sumir�?6OQ9ZO�O�O��?"F,3prens 8?�O�Ok_}_�"71_@C_�U_�_�_=�Kfurad/_�_U?�eowo
o�6�Csem?_recep�@8o�Jo�o�o�oo#6co��o�o�ocu� }�:�5drop�bdefeit�OIX���;8�z�t_1��I_�h�z���_23�E�W��������_3��ŏ׏h�z��_ �1�D�U������������Y͟^�p�������$SNPX_AS�G 2������� � 01%���Я � ?���PARAoM ����� �	��PӤr0Ө$�������OFT_KB_?CFG  ӣ�����OPIN_SI�M  ����}���������RVN�ORDY_DO � )�U���QS�TP_DSBi���ϐ�SR >�� � &#�D��O�O�:�TOP_?ON_ERRʿ��~o�PTN ������A��RING_PRMy��ܲVCNT_GP� 2��!���x 	����0��#���Gߔ�VD��RP 1��"�8Ѩ�*� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�}�z������� ��������
C@ Rdv����� �	*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?[?X?j?|?�?�? �?�?�?�?�?!OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLosopo �o�o�o�o�o�o�o  96HZl~� ������� ��2�D�V�`�PRG_�COUNTJ�眢�{�ENB��}�M���L���_UPD �1'�T  
 k������"�K�F�X� j���������۟֟� ��#��0�B�k�f�x� ��������ү����� �C�>�P�b������� ��ӿο����(� :�c�^�pςϫϦϸ� ������ ��;�6�H� Z߃�~ߐߢ������� ���� �2�[�V�h� z������������ 
�3�.�@�R�{�v��� ���������� *SN`r����t�_INFO 1=�Ҁ� 	 ��3�?��@������Z>����: B�J-���]��q9C�����'��f>>�` �AoB @{w �?�� >�@���9 �� DX��C���Z³��������YSDEBSUG����� dՉ��SP_PASSB?+LOG� ���  e� 9�  ���   UD1�:\;$�<"_MPACA-셽/�/����.쁝&SAV �D)��%d!|"�%��(SV�+TEM�_TIME 1�D'�� 0  Yq0���("�(��$&M7MEMBOK  �сd �d/�?�?�<X|NҀ� @�?v4�O :OJLOmOzI�J
! %@p1�O�O�O �O"3 __$_6_H_Z_l_ �n_�_�_�_�_@�_�_�_o"o\�e1o Vohozo�o�o�o�o�o �o�o
.@Rd`v���O5SK�0��8���?���F
ʉ1�H2OJ�A>J� ���u1h\O����(�O"�Oяb�ݏ��p�O�z0g� � ��0� f�x���~_K��Ο������$�C�7o g�y���������ӯ� ��	��-�?�Q�c�u�����������T1SVGUNSPD%%� '%��2M�ODE_LIM #a9"ܴ2�	�� D-۵ASK_?OPTION �9�!F�_DI ENB  U�%f��BC2_GRP 2!�u#o2��XB���C���ԼBCCF�G #��*< 8����`�@ I�4�Y��jߣߎ��� ����������E�0� i�T��x������� �����/��S�>�w�����t���u����� c���	B-f�. ��4[ ����� �� 02Dz h������� /
/@/./d/R/�/v/ �/�/�/�/�(���/? &?8?J?�/n?\?~?�? �?�?�?�?�?O�?4O "OXOFOhOjO|O�O�O �O�O�O�O__._T_ B_x_f_�_�_�_�_�_ �_�_oo>o�/Voho �o�o�o(o�o�o�o �o(:Lp^� ������� � 6�$�Z�H�~�l����� ��؏Ə��� ��0� 2�D�z�h���To��ȟ ���
���.��>�d� R�������z�Я���� ���(�*�<�r�`� ��������޿̿�� �8�&�\�Jπ�nϐ� �Ϥ������ϴ��(� F�X�j��ώ�|ߞ��� ���������0��T� B�x�f�������� ������>�,�N�t� b��������������� ��:(^�v� ���H���$ HZl:�~� ������2/ / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?P? R?d?�?�?�?t�?�? OO*O�?NO<O^O�O rO�O�O�O�O�O�O_ _8_&_H_J_\_�_�_ �_�_�_�_�_�_o4o "oXoFo|ojo�o�o�o �o�o�o�o�?6H fx���������v&��$TB�CSG_GRP �2$�u��  �&� 
 ?�  Q�c�M� ��q��������ˏ���*�1�&8�d�, �F�?&�	 �HCA�����b��CS�B�I�����V�>���ͪ�n�Ќ�ԝB���333��Bl"t������AÐ��fff:��.�C�����l�?�� ��G�w�R���A&��̧�����@��I�� -���
�X�u�@�R���轿̻�����	V�3.00I�	mt7���*� �%���ֶY��@f�f&� &�H�� �N� �O�  ������ ϏϘ�*�J2�1�'8��Ϥ�CFoG )�uB�Y E������d�9��#��#�I� W��pW�}�hߡߌ��� ���������
�C�.� g�R��v������ ��	���-��Q�<�u� `�r����������� I�cp"4��gR w������	 -?�cN�r ��&������ /</*/`/N/�/r/�/ �/�/�/�/?�/&?? J?8?Z?\?n?�?�?�? �?�?�?O�? OFO4O jOXO�O�O`�O�OtO �O_�O0__T_B_x_ f_�_�_�_�_�_�_�_ �_,ooPoboto�o@o �o�o�o�o�o�o�o( L:p^��� ����� �6�$� F�H�Z���~�����؏ Ə����2��OJ�\� n������������ ��
�@�R�d�v�4� ��������ί���� ү(�N�<�r�`����� ����ʿ̿޿��8� &�\�Jπ�nϐ϶Ϥ� ��������"��2�4� F�|�jߠߎ����߀� �� �߼�B�0�f�T� ��x��������� ���>�,�b�P����� ����v������� :(^L�p�� ��� �$H 6lZ|���� ��/�/ /2/h/ �߀/�/�/N/�/�/�/ 
?�/.??R?@?v?�? �?�?j?�?�?�?�?O *O<ONOOO�OrO�O �O�O�O�O�O _&__ J_8_n_\_�_�_�_�_ �_�_�_o�_4o"oXo Foho�o|o�o�o�o�o �o�/$6�/�ox f������� �,�>���t�b��� ����Ώ��򏬏�� &�(�:�p�^������� ��ܟʟ�� �6�$� Z�H�~�l�������د Ư��� ��D�2�T� z�h���Jȿڿ�� ����
�@�.�d�Rψ� vϬϾ����Ϡ���� ��*�`�r߄ߖ�P� �ߨ���������� &�\�J��n����� ��������"��F�4� j�X�z�|��������� ����0B�Zl ~(������ �,Pbt�D�������  9 # &0/�"�$TBJOP_GRP 2*���  �?�&	H"O#,vV,���� ן� =k% � Ȫ � �� ��$ @ g"	� �CA��&�?�SC��_%g!��"G��"k���/�+=�C�S�?��?��&0%0CR  B4��'??J7�/�/?33�3�2Y&0}?�:;���v 2�1�0-1*�20�6?�?20��7C�  D�!�,� �BL��OK:��Z�Bl  @pzB@�� s33C�1y �?gO  A�zG�2jG�&)A)E�O�J�;��|A?�f�f@U@�1C�Z0z8jO�Oz@���U�O��$fff0R)_;^;7xCsQ?ٶ4)@ �O�_tF�X_J\EU�_��V:�t-�Q(B� *@�Ooh�&-h$oZG Lo6oDoro�o~o8o�o �o�o�o3�oR@lVd��V4�&�`�q�%	V3.{00m#mt7A@��s*�l$!�'�� E��qE����E�]\E���HFP=F��{F*HfF@�D�FW�3Fp�?F�MF����F�MF���F�şF���F�=F����G�G�.8�CW�RD�3l)D��E�"��Ex�
E���E�,)F�dRFBFHF�n� F��F���MF�ɽF��,
GlG�g!G)�G�=��GS5�G�iĈ;��
;W�o�|& : E@Xz&/��&�"�?�0�&=;-E�STPARS  �(a E#HRw�A�BLE 1-V)� @�#R�7� (� �R�R�R�'T#!R�	R�
R�R�T��!R�R�R����RDI��`!���ԟ���
�r�O z���������̯ޮ��	Sx�^# <�����ÿ տ�����/�A�S� e�wωϛϭϿ����� ��;-w�{�_"��6�� 1�C�U���%�7�I��[����NUM  ��`!� �$  ��m���_CF�G .���!@�H IMEBF_T�T}���^#��G�VE�10m�H�]�G�R {1/�� 8��" �� �A�  ������������  �2�D�V�h�z����� ��������/
e @Rhv���� ���*<N `r������ '///]/8/J/`/n/@�/�/�/�/r���_���t�@~�t�MI_�CHANS� ~� ~!3DBGLVLS��~�s�$0ETHE�RAD ?��
w0�"��/�/�?�?�l�$0ROUTq��!�!�4�?�<SNMASKl8~�}1255.2E�s0O�BOTO�st�OOLO_FS_DI}��%�V9ORQCTRL� 0���#��MT �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo&l�OIo8omoq��PE_DETAI�J8�JPGL_CONFIG 6��ᄀ/cel�l/$CID$/grp1qo�o�o/壀�?Zl~ ���C����  �2��V�h�z����� ��?�Q����
��.� @�Ϗd�v��������� M������*�<�˟ ݟr���������̯@�}a���&�8�J�\���^o��c��`���˿ ݿ���Z�7�I�[� m�ϑ� ϵ������� ���!߰�E�W�i�{� �ߟ�.���������� ��A�S�e�w��� ��<���������+� ��O�a�s�������8� ������'9�� ]o����F� ��#5�Yk�}�����`��User Vi�ew �i}}12�34567890 �//,/>/P/X$� ,�cx/���2�U �/�/�/�/??s/�/�3�/b?t?�?�?�?�??�?�.4Q?O(O�:OLO^OpO�?�O�.5 O�O�O�O __$_�OE_�.6�O~_�_�_�_ �_�_7_�_�.7m_2o DoVohozo�o�_�o�.8!o�o�o
.@��oagr lCamera� �o����� �ޢE�*�<�N��h�z�`�������I  �v �)��$�6�H�Z�l� ���������؟���� �2�Y��vP9ɟ ~�������Ưد��� � �k�D�V�h�z��� ��E�W�I5�����  �2�D��h�zό�׿ ����������
߱�W� ދ��X�j�|ߎߠ߲� Y�������E��0�B� T�f�x�߁ulY��� ������
����@�R� d�������������� ��W� iy�.@Rd v�/����� *<N��W��i �������� /*/</�`/r/�/�/�/�/as9F/�/? ?1?C?U?�f?�?�? D/�?�?�?�?	OO-O
�j	�u0�?hOzO�O �O�O�Oi?�O�O
_�? ._@_R_d_v_�_/OAO �p�{,_�_�_oo)o ;o�O_oqo�o�_�o�o �o�o�o�_�u���o M_q���No� ��:�%�7�I�[� m�NEa����ˏݏ ����7�I�[��� �������ǟٟ���� ͻp�%�7�I�[�m�� &�����ǯ����� !�3�E�쟒�9�ܯ�� ����ǿٿ뿒��!� 3�~�W�i�{ύϟϱ� X�����H����!�3� E�W���{ߍߟ����������������  ��L�^�p���������� ��   "�*�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</�N/`/r/�/�  
���(  �@�( 	 �/�/�/�/ �/? ?6?$?F?H?Z?@�?~?�?�?�?�*2� �l�O/OAO�� eOwO�O�O�O�O��O �O�O_TO1_C_U_g_ y_�_�O�_�_�__�_ 	oo-o?oQo�_uo�o �o�_�o�o�o�o ^opoM_q�o�� ����6�%�7� ~[�m��������� ُ���D�!�3�E�W� i�{�ԏ��ß՟� ����/�A�S���w� ����⟿�ѯ���� �`�=�O�a������� ����Ϳ߿&�8��'� 9π�]�oρϓϥϷ� ��������F�#�5�G� Y�k�}��ϡ߳���� ������1�C�ߜ� y������������� 	��b�?�Q�c���� ����������(� )p�M_q������0@ �������� ��#�frh:\tpg�l\robots�\m10ia4_?7l.xml�X j|�������.��/1/C/U/ g/y/�/�/�/�/�/�/ �//?-???Q?c?u? �?�?�?�?�?�?�?
? O)O;OMO_OqO�O�O �O�O�O�O�OO _%_ 7_I_[_m__�_�_�_ �_�_�__�_!o3oEo Woio{o�o�o�o�o�o �o�_�o/ASe w�������o ��+�=�O�a�s����������͏ߏ��I �<<w  ?�� 4��,�N�|�b����� ��ʟ�Ο���0�� 8�f�L�~���������������(�$T�PGL_OUTP�UT 9����;� $�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ�����$�����2345678901��� � 2�D�V�^����υߗ� �߻�����w����'�9�K�]���}g��� ������o����1� C�U�g���u������� ����}���-?Q c������� ��);M_q 	������ �%/7/I/[/m/// �/�/�/�/�/�/�/? 3?E?W?i?{??%?�? �?�?�?�?O�?OAO SOeOwO�O!O�O�O�O��O�O_�O� $$Ӣ��OW=_o_ a_�_�_�_�_�_�_�_ �_#ooGo9oko]o�o �o�o�o�o�o�o�oC5g}��� �����}@���"�� ( 	 iW�E�{�i����� Ï��ӏՏ���A� /�e�S���w������� �џ���+��;�=��O���s����Ƹ  <<\ޯ� )�ͯ�)��M�_��� ʯ����<���ؿ��Ŀ � �~�$�V��Bό� ��x�����2ϼ�
ߤ� ��@�R�,�v߈���p� ����j�������<� �߬�r������ �����`�&�8���$� n�H�Z���������� ����"4Xj�� R��L���� |Tf �� v��0B//� &/P/*/</�/�/��/ �/h/�/??�/:?L? �/4?�??n?�?�?�? �? O^?�?6OHO�?lO ~OXO�O�OO$O�O�O �O_2___h_z_�O �_�_J_�_�_�_�_o�.o��)WGL1�.XML�cm�$�TPOFF_LI�M Š�p��{�qfN_SVy`�  �t�jP_�MON :����d�p�p2miS�TRTCHK �;���f~tbVT?COMPAT�h*q��fVWVAR �<�mMx�d R e�p�bua�_DEFPROG� %�i%C�OLOCA_ME�SA_IRVIS�I�`�rISPL�AY�`�n�rINST_MSK  �|� �zINUSsER �tLCK)���{QUICKMEx�pO��rSCREl����+rtpsc�t)������b���_��STz�iRA�CE_CFG U=�iMt�`	nt�
?��HNL C2>�z���T{ zr @�R�d�v����������К�ITEM 2�?,� �%$1�23456789y0�%�  =<�xC�U�]�  !c�k�wp'���ns�ѯ 5����k������j� ů��鯕���A�1�C� U�o�y�󿝿I�oρ� 忥�	��-ϧ�Q��� #�5ߙ�A߽�����e� �������M���q߃� L��g��ߋ���� %�w� �[���+�Q� c���o��������3� ��{�;������ G_����/�S e.�I�m� ��=�a/ 3/������k/ /�/�/�/]/?�/�/ �/?�/u?�?�??�? 5?G?Y?�?+O�?OOaO �?mO�?�?�OO�OCO __yO+_�O�Ox_�O �_�O�_�_�_?_�_c_ u_�_o�_Wo}o�o�_ �oo)o;o�o�oqo1 C�oO�o�o�� %��[��Z���S�@��_��g  ے_� ����y
 Ï�Џ����UD1:\����q�R_GR�P 1A �� 	 @�pe�w��a���������ߟ͞� ���ّ�>�)�b�M�?�  }���y� ����ӯ������	� �Q�?�u�c���������Ϳ�	-���~o�SCB 2B{� h�e�wωϛ���Ͽ�������e�UT�ORIAL C�{��@�j�V_CONFIG D{����������O�OUT?PUT E{����������� %�7�I�[�m���� �����������%� 7�I�[�m�������� ��������!3E Wi{������ ��/ASe w������� //+/=/O/a/s/�/ �/�/�/�/��/?? '?9?K?]?o?�?�?�? �?�?�/�?�?O#O5O GOYOkO}O�O�O�O�O �O�?�O__1_C_U_ g_y_�_�_�_�_�_�O �_	oo-o?oQocouo �o�o�o�o�o�_�o );M_q�� ����yߋ���� -�?�Q�c�u������� ��Ϗ���o�)�;� M�_�q���������˟ ݟ� ��%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���
� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� �1CUgy� ������	 -?Qcu��������/�x���$/6/ !/a/ ��/�/�/�/�/�/�/ ??'?9?K?]?�? �?�?�?�?�?�?�?O #O5OGOYOkO|?�O�O �O�O�O�O�O__1_ C_U_g_xO�_�_�_�_ �_�_�_	oo-o?oQo cot_�o�o�o�o�o�o �o);M_q �o������� �%�7�I�[�m�~�� ����Ǐُ����!� 3�E�W�i�z������� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�o�~���$TX_SCR�EEN 1F8%�  �}��~���������
�� ��m&��\�n߀ߒߤ� ��-�?������"�4� F��j��ߎ����� ����_����0�B�T� f�x����������� ����>��bt ����3�W (:L^��� �����e/� 6/H/Z/l/~/�//�/��$UALRM_�MSG ?����� �/���/�/)? ?M?@?q?d?v?�?�?��?�?�?�?O�%SEoV  �-EF��"ECFG Hv����  ���@�  AuA  w Bȁ�
 O ���ŨO�O�O�O�O_�_&_8_J_\_jWQAG�RP 2I[K 0��	 �O�_� �I_BBL_NO�TE J[JT?��l�����g@�RDEFP�RO� %�+ (�%SEGURA�_BAR"`REC_EPTOR�^%O VoAozoeo�o�o�o�o��o�o�o@�[F�KEYDATA �1K�ɞPp jG���_������z,(�����OINT  ]'�.)�DI+`TS�~��(INg���5�C�HOICEB���  TRINGS׏ ؏�'��K�2�o��� h�����ɟ۟����#�5��Y��y���/frh/gui�/whiteho?me.pngd���p��Ưدꯀ  |�point���0��B�T�f���{�direc�����ƿؿ4���{�in��#��5�G�Y�k�򯀡choic��ϰ������������strings�0�B�T�f�x�>��arwrgϲ� �������߉��)�;� M�_�q������� �������%�7�I�[� m������������� ����3EWi{ ������ �/ASew�� r������/!/ (E/W/i/{/�/�/./ �/�/�/�/??�//? S?e?w?�?�?�?<?�? �?�?OO+O�?OOaO sO�O�O�O8O�O�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5o�_Goko}o�o�o �o�oTo�o�o1 C�ogy���� P��	��-�?�Q� �u���������Ϗj�-܋�u�܏�@(�s��Q�c�r�,I����A�OINT  �]���� OOK �Tß�}�NDIR�ECܟ�  CH�OICE�����UCHUPG�H�s��� ~�����߯�د��� 9�K�2�o�V��������ɿ��whitehom����%�7�xI�X��poin����ϟϱ�����d�i/look}��(��:�L�^�i�indirec|Ϙߪ߼���|��g�choic����� �2�D�V�h�k�t?ouchup�ߠ���������g�arwrg��"�4�F�X�j� a�������������w� 0BTfx ������� ,>Pbt�� ����/�(/:/ L/^/p/�//�/�/�/ �/�/ ?׿�/6?H?Z? l?~?�?�/�?�?�?�? �?O�?2ODOVOhOzO �O�O-O�O�O�O�O
_ _�O@_R_d_v_�_�_ )_�_�_�_�_oo*o �_No`oro�o�o�o7o �o�o�o&�oJ \n����E� ���"�4��X�j� |�������A�֏��� ��0�B�яf�x��� ������O������h,�>�<L������u�����q���ͯ��,������ "�	�F�X�?�|�c��� ����ֿ������0� �T�f�Mϊ�qϮϕ� ���������,�>�? b�t߆ߘߪ߼�˟�� ����(�:�L���p� �������Y��� � �$�6�H���l�~��� ��������g���  2DV��z��� ��c�
.@ Rd������ �q//*/</N/`/ ��/�/�/�/�/�/�/ /?&?8?J?\?n?�/ �?�?�?�?�?�?{?O "O4OFOXOjO|OSߠO �O�O�O�O�OO_0_ B_T_f_x_�__�_�_ �_�_�_o�_,o>oPo boto�oo�o�o�o�o �o�o:L^p ��#���� � ��6�H�Z�l�~��� ��1�Ə؏���� � ��D�V�h�z�����-� ԟ���
��.��� R�d�v�������;�Я �����*���N�`�@r����������@�����@�������	��+�=��, )�n�!ߒ�y϶��ϯ� �����"�	�F�-�j� |�cߠ߇����߽��� ����B�T�;�x�_� ���O�������� ,�;�P�b�t������� ��K�����(: ��^p����G �� $6H� l~����U� �/ /2/D/�h/z/ �/�/�/�/�/c/�/
? ?.?@?R?�/v?�?�? �?�?�?_?�?OO*O <ONO`O�?�O�O�O�O �O�OmO__&_8_J_ \_�O�_�_�_�_�_�_ �_��o"o4oFoXojo q_�o�o�o�o�o�o�o �o0BTfx �������� ,�>�P�b�t������ ��Ώ������(�:� L�^�p��������ʟ ܟ� ����6�H�Z� l�~������Ưد� �����2�D�V�h�z� ����-�¿Կ���
� ϫ�@�R�d�vψϚ� )Ͼ���������*��`,��`���U�g�y�Qߛ��߇�,���ߑ���� &�8��\�C���y� ������������4� F�-�j�Q���u����� �������_BT fx������� �,�Pbt ���9���/ /(/�L/^/p/�/�/ �/�/G/�/�/ ??$? 6?�/Z?l?~?�?�?�? C?�?�?�?O O2ODO �?hOzO�O�O�O�OQO �O�O
__._@_�Od_ v_�_�_�_�_�___�_ oo*o<oNo�_ro�o �o�o�o�o[o�o &8J\3��� ����o��"�4� F�X�j��������ď ֏�w���0�B�T� f�����������ҟ� �����,�>�P�b�t� �������ί�򯁯 �(�:�L�^�p���� ����ʿܿ� Ϗ�$� 6�H�Z�l�~�Ϣϴ� ��������ߝ�2�D� V�h�zߌ�߰����� ����
��.�@�R�d��v���qp���>qp������� ��������,	N� r�Y����������� ����&J\C �g������ �"4X?|� m�����/� 0/B/T/f/x/�/�/+/ �/�/�/�/??�/>? P?b?t?�?�?'?�?�? �?�?OO(O�?LO^O pO�O�O�O5O�O�O�O  __$_�OH_Z_l_~_ �_�_�_C_�_�_�_o  o2o�_Vohozo�o�o �o?o�o�o�o
. @�odv���� M����*�<�� `�r���������̏� ����&�8�J�Q�n� ��������ȟڟi��� �"�4�F�X��|��� ����į֯e����� 0�B�T�f��������� ��ҿ�s���,�>� P�b��ϘϪϼ��� ���ρ��(�:�L�^� p��ϔߦ߸������� }��$�6�H�Z�l�~� ������������  �2�D�V�h�z�	��������������
�������5GY1{�g,y�q�� �<#`rY�} �����/&// J/1/n/U/�/�/�/�/ �/�/�/ݏ"?4?F?X? j?|?���?�?�?�?�? �?O�?0OBOTOfOxO �OO�O�O�O�O�O_ �O,_>_P_b_t_�_�_ '_�_�_�_�_oo�_ :oLo^opo�o�o#o�o �o�o�o $�oH Zl~��1�� ��� ��D�V�h� z�������?�ԏ��� 
��.���R�d�v��� ����;�П����� *�<�?`�r������� ����ޯ���&�8� J�ٯn���������ȿ W�����"�4�F�տ j�|ώϠϲ�����e� ����0�B�T���x� �ߜ߮�����a���� �,�>�P�b��߆�� �������o���(� :�L�^���������� ������}�$6H Zl������� �y 2DVh�zQ�|�Q�����������,�/./�/R/ 9/v/�/o/�/�/�/�/ �/?�/*?<?#?`?G? �?�?}?�?�?�?�?O O�?8OO\OnOM��O �O�O�O�O�O�_"_ 4_F_X_j_|__�_�_ �_�_�_�_�_o0oBo Tofoxoo�o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� ��#���ʏ܏� �� ��6�H�Z�l�~���� ��Ɵ؟���� ��� D�V�h�z�����-�¯ ԯ���
����@�R� d�v��������Oп� ����*�1�N�`�r� �ϖϨϺ�I������ �&�8���\�n߀ߒ� �߶�E��������"� 4�F���j�|���� ��S�������0�B� ��f�x����������� a���,>P�� t�����]� (:L^�� �����k // $/6/H/Z/�~/�/�/��/�/�/�/���+}������?@'?9=?[?m?G6,YO �?QO�?�?�?�?�?O O@ORO9OvO]O�O�O �O�O�O�O_�O*__ N_5_r_�_k_�_�_�_ �_��oo&o8oJo\o k/�o�o�o�o�o�o�o {o"4FXj�o ������w� �0�B�T�f�x���� ����ҏ������,� >�P�b�t�������� Ο������(�:�L� ^�p��������ʯܯ � ���$�6�H�Z�l� ~������ƿؿ��� ϝ�2�D�V�h�zό� ϰ���������
�� �_@�R�d�v߈ߚߡ� ����������*�� N�`�r����7��� ������&���J�\� n���������E����� ��"4��Xj| ���A��� 0B�fx�� ��O��//,/ >/�b/t/�/�/�/�/ �/]/�/??(?:?L? �/p?�?�?�?�?�?Y?��? OO$O6OHOZO��$UI_INUS�ER  ����{A� � [O_O_ME�NHIST 1L�{E  �( �@��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1`�O__1_C_�'�O��N71�@BARR�A_ESTEIRAA�O�_�_�_�39X_��Eedit�BCO�LOCA�@SA_�IRVISION �_$o6oHo�1)�_�O527o�o�o�o�o]ooo�d2�o0B��o� �o�m936 �o����dv�A48#�5�G�Y�����O����ŏ׏�5���0�A����"�4� F�X�j�m��������� ȟڟ�{��"�4�F� X�j���������į֯ �w���0�B�T�f� x��������ҿ��� ���,�>�P�b�t�� �Ϫϼ��������� (�:�L�^�p߂߅�#� �������� ���6� H�Z�l�~������ ����������D�V� h�z�����-������� ��
��@Rdv ��);��� *�N`r�� �����//&/ 8/�\/n/�/�/�/�/ E/�/�/�/?"?4?F? �/j?|?�?�?�?�?S? �?�?OO0OBO�?fO xO�O�O�O�O�OaO�O __,_>_P_;t_�_ �_�_�_�_�_�Ooo (o:oLo^o�_�o�o�o �o�o�oko $6 HZl�o���� ��y� �2�D�V� h��������ԏ� �����.�@�R�d�v��aX�$UI_PA�NEDATA 1�N������  	�}�1/frh/vi�sion/vsv�trn.stm?�_screen_�id=2&_fo�cus_flag�=1 =TP&_�lines=15�&_column�s=40ڑnt=�24&_page�=wholede�v��\V)pri9m#�L�  }O�s�`��������ͯ )ϯ �گ���;�M�4�q� X�������˿������%�\V�� �    �f]���cgt?p/flex�ɓ�width=�h�eight=10��ice�ِ��3���1
�dou�b�2/��ual ����_��"�4�F�X� j�ώ�u߲��߫��� �����B�)�f�M�����3� D�?  ����� ��*�<�N�`���� �Ϩ���������i� &8\C��y ������4Xj������� ����� /S$/ ��H/Z/l/~/�/�/	/ �/�/�/�/�/ ?2?? V?=?z?a?�?�?�?�? �?�?
O}�@OROdO vO�O�O�?�O1/�O�O __*_<_N_�Or_Y_ �_}_�_�_�_�_�_o &ooJo1ono�ogo�o O)O�o�o�o"4 �oXj�O���� ��O��0�B�)� f�M������������ ��ݏ��>��o�o� ��������Ο��3�� w(�:�L�^�p���� ������ܯï ���� 6��Z�A�~���w��� ��ؿ�]�o� �2�D� V�h�z�Ϳ������� ����
��.ߕ�R�9� v�]ߚ߬ߓ��߷��� ���*��N�`�G����	�������������"�)��G���6�s� ����������4����� ��K2oV� �������#������$UI_�POSTYPE � ��� 	 /�UQ�UICKMEN � ds�WR�ESTORE 1�O�  O��� /#���m+/T/f/x/ �/�/?/�/�/�/�/? �/,?>?P?b?t?/�? �?�??�?�?OO(O �?LO^OpO�O�O�OIO �O�O�O __�?_1_ C_�O~_�_�_�_�_i_ �_�_o o2o�_Voho zo�o�oI_So�o�oAo �o.@Rd� ����s��� *�<��oI�[�m���� ��̏ޏ�����&�8� J�\�n��������ȟ�ڟ�SCRE�?��u1s]c�u2�3�U4�5�6�7��8��TAT`�� ��MUSE1R�����ks���U3��4��5��6���7��8��UNDO_CFG PdX����UPDX�����None����_INFO �1Q�<��0%��W���E���i��� ������տ���:� L�/�pς�eϦύ)��OFFSET 	Td@���{���� ��	��-�Z�Q�cߐ� �ߙ��ϝ������� � �)�V�M�_�q�۹�����
���t���)�WORK U4�����A�S��ψ��UFRAME  ����&�RTOL_ABRT��$����ENB����GRP� 1V��Cz  A��� +=Oas�����U������MSKG  �<���N��%4��%��)��O_EVN������>�2W��
 h���UEV��!�td:\eve�nt_user\�-�C7���}�F���SP��spotweld�!C6����!�Z/�/:'� H/~/l/�/�/�/�/-? �/Q?�/? ?�?D?�? h?z?�?O�?)O�?�? OqO`O�O@ORO�OvO �O_�O�O7_�O[__4Z]W+�2X����#8V_�_�_ �_�_ o�_,o>oobotoOo �o�o�o�o�o�o �o:L'p�]�����$VARS�_CONFI�Yn�� FP{���|oCCRG�\�ʨ>�{�t�D� �BH� pk�a�C�2� ��}�?���C,�&Q=��ͩ�A ��MR2b����	}�	��@�%�1: SC13?0EF2 *�����{�����X� �5�}�����A@k�C��F� w�Q� [���|����������"T����\�ϟ ��\� B��� ;�e�@�ǟ`�����S� ����̯���ۯ�&� }��\�G�Y���E���\ȿ�TCC�c
Е�������pGFt�pgd��-��23456789�017�?��ׁ$���4�v�Nm�� ��ς��BW�����i�}�:�o=LA�څ� 6�@�6�ͿZ���i�7�	���(��W���-�]� X�jĈߚߕϳϹ��� ������%�7�I�r� m�ߨ�ߵ������� ���8�3�E�W���� ��}��������������/�A�S�e�w��MgODE��t �RSLT e�|k�%"zς��;��1��d��`��S�ELEC��c���	IA_WO�Puf �� W,		������G�P ������RTSYNCSE� ��$�	#WIN?URL ?*ـ�;\/n/�/�/�/��/�uISIONT�MOU���A# ���%�gSۣ��SۥP�� �FR:\�#\DA�TA\�/ ��� MC6LOG�?   UD1�6EX@?\�' B@ ���2�T1  abriel_Fariak?�P5�?�?����� �n6  ���xGV�2\� -��5>��   ��Z��@U058TRAI�Nj?��*B{Rd_C�p��D #`�{2��'$�"��h#� (�kI�Mw��O�O �O�O�O1__U_C_]_�g_y_�_�_�_�(STA� i��@�o o�2oI8$>obo�%_G�E�j#��~@ ��
�\��btgHO�MIN�kSۮ���`�2,,��C�WǖBveJMPE�RR 2l#�
  ��I:��"�4 Fwj|����������&%S_�g0RE�m�^۴L�EXdn�1-�ehoVMPHASOE  �e׃B�ޱOFF _EN�B  �$VP}2�$oSۯ��)x�c C;�@ �ax;���?s33'D*AA��]� ��(0ޱ�`r}�XC���܅��� ��[��6�������6��]���>�VYD-۟E �B�[�t\1�6��+FV����W��5 d�����,�>�'Es����W�I�ǟ���  ��I�����9�k�ɯ ;�������ׯɿ3�տ ����C�8�g�Yϋ��� ����ϱϿ�����-� "�Q�c�u�jߙ�?��� �ߩ߻����u���M� B�T��u��߁��� ������7�,�[�m� ��]�k�}��������� �!�E�����CU g���!����  /!�-WQ�� ����c	/�/)/?/M's�TD__FILTE�`s�kg �x2�`��� �/�/�/�/�/	??-? ??Q?�6�/~?�?�?�?��?�?�?�?O OoiS�HIFTMENU� 1t}<5�% 5�~O)�\O�O�O�O�O �O�O�O'_�O_6_o_�F_X_�_|_�_�_�_�	LIVE/SN�AP�Svsflsiv���_�z`/ION ҀU
`bmenu&o+o�_�oP�oV"<E�uz��4IkMO�v���zq��WAITDINEND  �ec��b��fOKوOUT��hSDyTIM.du��o|G�} #�{C�zb�z�x�RELE��ڋxT�M�{�d��c_A�CT`و��x_D?ATA wz����%  EGA_T�ORNO�o.Mx�R�DIS
`E��$�XVR�ax�n��$ZABC_GRoP 1yz���� ,�2̏.MZ�D��CSCH�`zd���aP@�h@�IP�b{'����şן�[�MPCF__G 1|'���A0�r�8��� �}'��(�p�s� 	|(���  <l0�  4�13c�c�?�  ��5� )o��3��ﲯ��cc��� DX���C��Z�>w�?��}�*�����@(������,&��� ����ɯۯ������o���w���� /�³��۰�c̿޷ĸ���	��1�@?�i���'�9�0?��Q��	��`~����_�CYLIND~!�� Р ,(  *.�?ݧ+�0h�Oߌ�s� ���� ����(�	�x�-��&� c�߇�������j� P����)��~�_�q���� �2�'��� �&�����������&��I��cA����SPHERE 2������� ���A�T/A�� e����� �/N`=/�a/H/�Z/�/��/�/�/��Z:�� ��f