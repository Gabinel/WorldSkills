��   g�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����BIN_CFG_�TX 	$EN�TRIES  �$Q0FP?N�G1F1O2F2�OPz ?CNET�G���DHCP�_CTRL. � 0 7 ABL�E? $IPUS~�RETRAT��$SETHOS�T��NSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM�� !� FT�� @� LOG_�8	,CMO>$�DNLD_FIL�TER�SUBDIRCAPC��\8 . 4� H�{ADDRTYPz�H NGTH�̉��z +LS�q D $R�OBOTIG �P�EER�� MAS�K�MRU~OM�GDEV��PI�NFO�  {$$$TI ��RCM+T A$( </�QSIZ�!�S� TATUS_�%$MAILSE�RV $PLA�N� <$LIN><$CLU���<$TO�P$C�C�&FR�&YJE�C|!Z%ENB �� ALAR:!BF�TP,�#,V8 }S��$VAR�)�M�ON�&���&A7PPL�&PA� �%���'POR�Y#_|�!�"ALERT�&�i2URL }>Z3ATTAC��0�ERR_THRO�U3US�9H!�8� CqH- c%�4MAX?wWS_|1��1'MOD��1I�  ��1o (�1PWD  � LA��0��ND�1TRYFD�ELA-C�0G'AE�RSI��1Q'RO.BICLK_HM 0Q'ί XML+ 3SG�FRMU3T� !O�UU3 G_�-COAP1�F33�AQ'C[2�%�B_AU�� 9 �R�!UPDb&P�COU{!�CFO 2 
$V*W8�@c%ACC_HYQ�SNA�UMMY�1oW2"$DM*�  $DIS��SM	 !l5�o!�"%Q7�IDZP�%� �VR�0z�UP� _DLVS�PAR�  �S)N,#
3 �_�R�!_WI�CTZ_�INDE�3^`OFYF� ~URmiD��)c�   ts Z!`MON�r�cD��bHOUU#�E%A�f�a�f�a�fL�OCA� #$N�S0H_HE��r�@I�/  d8`�ARPH&�_IP�F�W_* O�F``QFAsD90�V�HO_� 5R42PS�Wq?�TEL�# P���90WWORAXQE� �LV�[R2�IcCE��p� �$cs  ����qJ��
��
�p�PS�A��w# 0�	�Iz0AL��'� �
���F��p��!�p�i��$� 2Q�$a���@������ Q���!�q�����$� _FL�TR  �\� U�����������$Q�2��7rSH^`D 1Q� P㏙�f���ş�� 韬��П1���=�� f���N���r�ӯ���� ���ޯ�Q��u�8� ��\�������󿶿� ڿ;���_�"�Xϕτ� ��|��Ϡ������� 6�[���Bߣ�f��� ���߮���!���E�� i�,��P�b������ �����/���(�e�T�`��L�����z _LUA�1�x!1."��0��p���1��p�255.0��r��n���2����d  %7I[3e��@� ����[4����T'9[5 U���{���[6���D �//)/�s��QȁMA���MA� ������ Q� ��u.<�/?&? �/J?\?n?A?�?�?m�P�?�?�?�?�?O.O�@OROOvO�O�Ou.�kOl�q��O�L
Z�DT Statu�sZO�O5_G_Y_n�}�iRConnect: irc{T//alert^ �_�_�_�_mW#_oo�,o>oPobot�^�d~2g���go�o�o�o �o�o�o	-?Q�cul�$$c96�2b37a-1a�c0-eb2a-�f1c7-8c6�eb584036�`(�_�_����"�p�1!W��(� �"S��JE�� X��C� ��,$���W��� ˏ���֏��%��I� 0�m��f�����ǟ��@�����!��u�R�s���� DM_�!�����SMTP�_CTRL 	����%����DF� ��ۯt�ʯ��'��Lz�N��!
j��y��q�u���������#L�USTOM' j������ � ���$TCPIPd�j��H�%�"��EL�����!�>��H!TP��j��rj3_tp��b;���i�!K�CLG�L�i���5�!CRT�ϔ����"�u�!CONS���M�[�ib_s'mon����