��   K�A��*SYST�EM*��V9.3�044 1/9�/2020 A� 	  ����CELL_GRP�_T   � �$'FRAME� $MOU�NT_LOCCC�F_METHOD�  $CPY�_SRC_IDX�_PLATFRM�_OFSCtDI�M_ $BASE{ FSETC���AUX_ORDER   ��XYZ_MAP ��� �LE�NGTH�TTC?H_GP_M~ a �AUTORAIL�_���$$CL�ASS  �S����D��DVERSION�  0��/IRTUAL�-9LOOR qG��DD<x$?������k, � 1 <DwX�< y�����C������	/�� Z�Zm//�/_/�/8�/�/$ �/�/|	?';�$MNU>YA\"�  <����;8_���4�g0U���߶X��k0�5�;�s0�D	}�����àW���0�?/�?'�? �?�?�?�?!OO)OWO =OOO�OsO�O�O�O�O �O_�O_A_'_�;5�NUM  ���x�w92TOOLC?\ 
Y8&/V_��B45_�_o/_o=o #o5oWo�oko�o�o�o �o�o�o�o9A oU������ qX�Q�Vy�[