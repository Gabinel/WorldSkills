��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@��&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	4SU�SRVI 1  < `�R*�R�n�QPRI�m� �t1�PTRIP�"m��$$CLASP ����a��R2��R `\ SI�	g�  0�aIRTs1	o`�'2 L1�L1���R	 ,��?���a1`��b�ba ����� � y�o��
 ��a��o�o1CU  �oz�����c �
��.�@�R��v� ��������Џ�q�� �*�<�N�`���� ����̟ޟm���&� 8�J�\�n��������� ȯگ�{��"�4�F� X�j���������Ŀֿ����`TPTX�����/�`� sȄ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ��� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F�X���|��������������a�f�b�� ($p�-����T�?�x���a�a��c���c����l��c�g���aR�ah�ah��at2�h�	f�����������`���` � ���f epS��h#h�F�brc Xc�B 1)h�R \ _��� RE�G VED]����wholemod�.htm�	sin�gl	doub~ trip8browsQ �����u�� �//@/���_dev.sl�/43� 1�,	t�/_ �/;/i/??/?�/S?�e?w?�?�?�?�  ��?�?OO%O7OIO0[OmOO�E @�?�O �O�O�O�O_�F�	�? �?;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omooM'�o�o�o �o�o�o+=O as������ ���?>�P�b�t��� ������Ώ���O�� ���L�^�_'_��� ����ş�����6� 1�C�U�~�y�����Ư ��ӯ�o���-�?� Q�c�u���������Ͽ ����)�;�M�_� -��ϬϾ�������� �*�<�7�`�r�A�S� �ߺ�q���i����� !�J�E�W�i���� ����������"��/� ��O�I�w��������� ������+=O as������� ,>Pbt� ��߼���// �����^/Y/k/}/�/ �/�/�/�/�/�/?6? 1?C?U?~?y?�?Y��? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__�R_d_v_ �_�_�_�_�_�_�_��o*o�_o`oro�j��$UI_TOPMENU 1K`��aR 
�d�a*Q)*d?efault5_]�*level�0 * [	 ��o�0�o'rtpio[23]�8tpst[1[x�)w9�o	�=h�58E01_l.�png��6me�nu5�y�p�13�z��z	�4���q��]���������̏ ޏ)Rr���+�=�O��a���prim=��page,1422,1h�����ş ן����1�C�U��g���|�class,5p�����ɯۯ4�����13��*��<�N�`�r���|�53������ҿ�����|�8��1�C�U�g� y����ϯ���������"Y�`�a�o/��m!�`�q�Y��avtyl}<Tfqmf[0nl�}	��c[164[w��59[x�qG�y��tC8�|�29��o� %�1���{��m��!� ����0�B���f�x����������o���80 ��'9K~���2P�����\ ��'9K�� ����������1��/$/6/H/Z/U��|�ainedi�'ߑ/�/�/�/�/P��config=s�ingle&|�wintp���/$?6?�H?Z?	�ߐ??ٷ�gl[57�ٳq��?H�;gp�08�ݲ07I��?F��F2JO[6��:�?)O�O�x �� �4s�x�O��� $��`�o�H_Z_l_~_ �_�_Q��_�_�_�_o  o�_DoVohozo�o�o��o�!;�$doub�5o��13��&d�ual�i38��,!4�o&�o9�o�n �o�a8���Ao�@���&�8��%3L!=}!��o�b8@��� ������z���(��:��+:T��i48,�2o��b{����ʟ {?�;�M�sc���;���s�� �}���e�au��X��@�F7L���`�O��2�h�z�6e�u7�����ｿϿ`���̏�27�� G�Y�k�}Ϗ��0�s@���������!�1�M�_�q߃ߕ�� �����������7� I�[�m��������������!�����6 (�]�o��������$��746�����)��C�ߟT�	TP?TX[209�<A�w2IHJ���Bw1 H�]H�����02��A#��[Ttv`��O�L#_��0� \��5S[�tr?eeview3v��3��~�381,26M/_/q/0�/�/ �/�/�/�/~/?%?7? I?[?m?�o/(��o5%0���?�?�?�A�?\1~��?8"2��eOwO �?�?(}�LEK��O�O _�O��8@�ONOa_s_�_��6_d�E_�_�_ �_oV�#_���_�So oo�o�oB�o�o��o A�oq+=O as��o���� ���(�9���Q�x� ��������ҏ?��� �,�>�P�ߏt����� ����Ο]�����(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z��l�������ƿؿ �y�� �2�D�V�h� ���Ϟϰ������ϕo �o��o@ߧE�c�u� �ߙ߽߬�����O��� �)�<�M�_�q��� W���������&�8� ��\�n���������E� ������"4��X j|����S� �0B�fx ����O��/ /,/>/P/�t/�/�/ �/�/�/]/�/??(? :?L?��߂?1ߦ?� ���?�?�?�?O$O5O GO�?SO}O�O�O�O�O �O�O�O��2_D_V_h_ z_�_�_�/�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� 7�����&�� J�\�n���������E� ڏ����"�4�ÏX� j�|�������a?s?� �?�sO_/�A�S�e� w������������� ��,�=�O�a�#_�� ����ο��=��(� :�L�^�pς�Ϧϸ� ������ ߏ�$�6�H� Z�l�~�ߐߴ����� ������2�D�V�h� z������������ 
����@�R�d�v��� ��)����������ƚԔ*defa�ult%��*level8�ٯw����? tp�st[1]�	�y��tpio[23���u����J\menu7�_l.png_&|13��5�{4�y4�u6��� //'/9/K/]/���/ �/�/�/�/�/j/�/?�#?5?G?Y?k?�"p�rim=|pag?e,74,1p?�?��?�?�?�?�"�6class,13�?�*O<ONO`OrOOB5�xO�O�O�O�O�O�# L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]o�oo�o`�$UI_�USERVIEW� 1֑֑�R 
�� �o��o�o[m�o '9K] ��� ��l���#�5� �oB�T�f������ŏ ׏鏌���1�C�U� g�
���������ӟ~� ����v�?�Q�c�u� ��*�����ϯ�󯖯 �)�;�M�_�
��~� �����ݿ���%� ȿI�[�m�ϑ�4ϵ� �������Ϩ�
��.� ��i�{ߍߟ߱�T��� ������/���S�e� w���Fߨ����>� ��+�=�O���s��� ������^����� '����FX��|� �����#5 GY�}���� p���h1/C/U/ g/y//�/�/�/�/�/ �/�/?-???Q?c?/ p?�?�??�?�?�?O O�?;OMO_OqO�O&O �O�O�O�O�O�?�O_  _�OD_m__�_�_�_ X_�_�_�_o!o�_Eo Woio{o�o0h