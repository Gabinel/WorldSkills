��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@��&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	4SU�SRVI 1  < `�R*�R�n�QPRI�m� �t1�PTRIP�"m��$$CLASP ����a��R2��R `\ SI�	g�  0�aIRTs1	o`�'2 L1�L1���R	 ,��?���a1`��b�d~a���� � �`y�o��
 ��a��o�o1CU  �oz�����c �
��.�@�R��v� ��������Џ�q�� �*�<�N�`���� ����̟ޟm���&� 8�J�\�n��������� ȯگ�{��"�4�F� X�j���������Ŀֿ����`TPTX�����/�`� sȄ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ��� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F�X���|��������������a�f�b�� ($p�-����T�?�x���a�a��c���c����l��c�g���aR�ah�ah��at2�h�	f�����������a���`  ����f ep)��h#h�F�bc� Xc�B 1)hR_ \ _�� REG �VED]���w�holemod.�htm�	sing}l	doub �trip8?browsQ� ����u����//@/���d/ev.sl�/3� 1�,	t�/_�/ ;/i/??/?�/S?e?pw?�?�?�?� � �?�?OO%O7OIO[OmOO�E @�?�O�O �O�O�O_�F�	�?�? ;_M___q_�_�_�_�_ �_�_�_oo%o7oIo [omooM'�o�o�o�o �o�o+=Oa s������� ��?>�P�b�t����� ����Ώ���O��� ��L�^�_'_����� ��ş�����6�1� C�U�~�y�����Ư�� ӯ�o���-�?�Q� c�u���������Ͽ� ���)�;�M�_�-� �ϬϾ��������� *�<�7�`�r�A�Sߨ� ��q���i�����!� J�E�W�i����� ��������"��/��� O�I�w����������� ����+=Oa s������� ,>Pbt�� �߼���//�� ���^/Y/k/}/�/�/ �/�/�/�/�/?6?1? C?U?~?y?�?Y��?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__�R_d_v_�_ �_�_�_�_�_�_�o�*o�_o`oro�j�$�UI_TOPME?NU 1K`�a�R 
�d�a*Q)*de�fault5_]�*level0{ * [	 �o��0�o'rtp�io[23]�8?tpst[1[x)�w9�o	�=h5�8E01_l.p�ng��6mencu5�y�p�13�z���z	�4���q��]���������̏ޏ )Rr���+�=�O�a�~��prim=��page,1422,1h�����şן ����1�C�U�g����|�class,5p�����ɯۯ�����13��*�<��N�`�r���|�53�������ҿ�����|�8��1�C�U�g�y� ���ϯ���������"Y�`�a�o/��m!ηq0�Y��avtyl}T�fqmf[0nl�	>��c[164[w�Ճ59[x�qG�y��tC	8�|�29��o�%� 1���{��m��!��� ��0�B���f�x���`������o���80��'9K~���2 P�����\�� '9K�������������1���/$/6/H/Z/U�~|�ainedi'���/�/�/�/�/P�c�onfig=si�ngle&|�wintp���/$?6?H? Z?!Z�a�h?�?�e�? ���?�?�?OO+O =OOO�?[O�O�O�O�O �O�O�O_a�%_L_^_ p_�_�_�_U��_�_�_  oo$o�_HoZolo~o �o�o1o�o�o�o�o  2�oVhz�� �?���
��.� �@�d�v��������� M�����*�<�ˏ�`�r���������^ ��;�M�sc���;����s�� �}���e�u0��X��@�F7L����`��t꒯4�j�X�6e�u7�����ｿϿ`������27�� G�Y�k�}Ϗ��0�s@���������!�1�M�_�q߃ߕ�T� �����������7� I�[�m��������������!�����6 (�]�o��������$��746�����)�t<ϯ\�5	TPTX[209©|Dw�24§J��
�w18��� ����02��A#��[	�tv`�RxL�u10�1���5S�:�$treevi�ew3��3��&d�ual=o'81,26,4�O/a/ s/2�/�/�/�/�/�/ �/?'?9?K?]?o?��	;/&�3$/6$���? �?�?
?#O5OGOYOkO�}O�?�? "2�?8"2@K��O�O_�O��1�?`�E��g_y_�_�6_��edit��>_P_ �_�_o��/���_�C ooo�o�oB�o�o� �oA�o�+= Oas��o��� ����(�9���Q� x���������ҏO�� ��,�>�P�ߏt��� ������Ο]����� (�:�L�^�ퟂ����� ��ʯܯk� ��$�6� H�Z��l�������ƿ ؿ�y�� �2�D�V� h����Ϟϰ������� �o�o��o@ߧE�c� u߇ߙ߽߬�����O� ���)�<�M�_�q�� ��W���������&� 8���\�n��������� E�������"4�� Xj|����S ��0B�f x����O�� //,/>/P/�t/�/ �/�/�/�/]/�/?? (?:?L?��߂?1ߦ? ���?�?�?�?O$O 5OGO�?SO}O�O�O�O �O�O�O�O��2_D_V_ h_z_�_�_�/�_�_�_ �_
oo�_@oRodovo �o�o)o�o�o�o�o *�oN`r�� �7�����&� �J�\�n��������� E�ڏ����"�4�Ï X�j�|�������a?s? 蟗?�sO_/�A�S� e�w����������� ����,�=�O�a�#_ ������ο��=�� (�:�L�^�pς�Ϧ� �������� ߏ�$�6� H�Z�l�~�ߐߴ��� ��������2�D�V� h�z���������� ��
����@�R�d�v� ����)����������ƚԔ*def�ault%��*?level8�ٯ�w���? t?pst[1]�	��y�tpio[#23���u����J\menu7_l.png_M|13��5�h{�y4�u6� ��//'/9/K/]/�� �/�/�/�/�/�/j/�/�?#?5?G?Y?k?�"�prim=|page,74,1p?@�?�?�?�?�?�"�6�class,13 �?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo�]ooo�o`�$UI�_USERVIE�W 1֑֑�R 
�A��o��o�o[m�o '9K] �� ���l���#� 5��oB�T�f������ ŏ׏鏌���1�C� U�g�
���������ӟ ~�����v�?�Q�c� u���*�����ϯ�� ���)�;�M�_�
�� ~������ݿ��� %�ȿI�[�m�ϑ�4� ���������Ϩ�
�� .ߠ�i�{ߍߟ߱�T� ��������/���S� e�w���Fߨ���� >���+�=�O���s� ��������^����� '����FX��| ������# 5GY�}��� �p���h1/C/ U/g/y//�/�/�/�/ �/�/�/?-???Q?c? /p?�?�??�?�?�? OO�?;OMO_OqO�O &O�O�O�O�O�O�?�O _ _�OD_m__�_�_ �_X_�_�_�_o!o�_ EoWoio{o�o0h