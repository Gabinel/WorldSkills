��   8��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_IOC�_T   P �$OPERAT�ION  $�L_TYPBID�XBR1H[ S2�]2R��$$C�LASS  �������P��P�� VERS?��  0�~�IRTUAL�ܡ' 2 �P @ ��  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt����������_C_C�CL ?�� � 	All �param��
�Base!�P�os./Speed checkF��Safe I/O� connect�}R��,�>�P�b�t�SI��@���� �,�>�g�b�t��� ������Ο����� ?�:�L�^��������� ϯʯܯ���$�6� _�Z�l�~�������ƿ �����7�2�D�V� �zόϞ��������� �
��.�W�R�d�v� �ߚ߬߾�������� /�*�<�N�w�r���@����������O� ���C�l�g�y����� ����������	D ?Qc����� ���);d _q������ �//</7/I/[/�/ /�/�/�/�/�/�/? ?!?3?\?W?i?{?�? �?�?�?�?�?�?O4O /OAOSO|OwO�O�O�O@�O�O�O__�}N�  7�_b_�_�_�_ �_�_�_�_�_oo(o :oco^opo�o�o�o�o �o�o�o ;6H Z�~��������� �+_�SI ��6�7���������ȏ �����9�4�F�X� ��|�����ɟğ֟� ���0�Y�T�f�x� ������������� 1�,�>�P�y�t����� ����ο�	���(� Q�L�^�pϙϔϦϸ� ������ �)�$�6�H� q�l�~ߐ߹ߴ����߀���� �I�D�O�P�C_�u�SFDII1N��2���3��4���5���6$���7���8-�`� Q�c�u����������� ����);M_ q������� %7I[m �������/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ ����)�;�M�_� q���������˟ݟ� ��%�7�I�[�f�x�	O���O�ﵣ�ﵣ �ﵣ�ﵣ�ﵣ��� ,���D�~�o������� ��ɿ�����:�5� G�Yς�}Ϗϡ����� �������1�Z�U� g�yߢߝ߯������� ��	�2�-�?�Q�z�u� ����������
�� �)�R�M�_�q����� ����������*% 7Irm��� ���!JE Wi������ ��"////A/j/e/ w/�/�/�/�/�/�/�/ ??B?=?O?a?�?�? �?�?�?�?�?�?OO 'O9ObO]OoO�O�O�O �O�O�O�O�O_:_5_ G_Y_�_}_�_�_�_�_ �_�_ooo1oZoUo�goyo�o��SI��޳�VOFF�oF�ENCE�oEX�EMG�o�osN�TED"OP�2qAUTO:�T��ysӯqM�CC�3pCSBP��
POSSP�D_ENBzC�ONF_OK�~F�_IPAR_CR(�z�g�������oB�q_�oY�pE��DIS�|C_D6�r_~��� 