��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@��&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	4SU�SRVI 1  < `�R*�R�n�QPRI�m� �t1�PTRIP�"m��$$CLASP ����a��R2��R `\ SI�	g�  0�aIRTs1	o`�'2 L1�L1���R	 ,��I?���b1`�c�c~a��  � �  <�o��
 ��a�o@�o1CU �o z�����c� 
��.�@�R��v��� ������Џ�q��� *�<�N�`������ ��̟ޟm���&�8� J�\�n���������ȯ گ�{��"�4�F�X� j���������Ŀֿ����`TPT�X�����/�`� sȄ�$/s�oftpart/�genlink?�help=/md�/tpmenu.dg���ϨϺ��υ� ����&�8�J���n� �ߒߤ߶���W����� �"�4�F�X���|��`����������ae�f�oC ($p�-����T�?�x��� a�a��oŪ����l��c�g���a�ah��h��a2�h�]	f�����������`���`  ����f ep���h#h�F�bc �Xc�B 1)hR� \ _��� REG V�ED]���wh�olemod.h�tm�	singl�	doub �trip8browsQ�� ���u���/�/@/���dev.sl�/3� 1�,	t�/_�/;/ i/??/?�/S?e?w?8�?�?�?� ��? �?OO%O7OIO[OmOO�E @�?�O�O�O �O�O_�F�	�?�?;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o mooM'�o�o�o�o�o �o+=Oas �������� �?>�P�b�t������� ��Ώ���O����� L�^�_'_������� ş�����6�1�C� U�~�y�����Ư��ӯ �o���-�?�Q�c� u���������Ͽ�� ��)�;�M�_�-��� �Ͼ���������*� <�7�`�r�A�Sߨߺ� q���i�����!�J� E�W�i������� ������"��/���O� I�w������������� ��+=Oas ������� ,>Pbt���� ����//���� �^/Y/k/}/�/�/�/ �/�/�/�/?6?1?C? U?~?y?�?Y��?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __�R_d_v_�_�_ �_�_�_�_�_�o*o��_o`oro�j�$U�I_TOPMEN�U 1K`�a�R 
d��a*Q)*def�ault5_]�*level0 =* [	 �o�0��o'rtpi�o[23]�8tpst[1[x)w�9�o	�=h58�E01_l.pn�g��6menu15�y�p�13�z���z	�4���q�� ]���������̏ޏ)R r���+�=�O�a����prim=�p�age,1422,1h�����şן� ���1�C�U�g����|�class,5p�����ɯۯ�����13��*�<�N�h`�r���|�53��@����ҿ�����|�8��1�C�U�g�y�����ϯ���������"Y �`�a�o/��m!ηq�Y��avtyl}TfqOmf[0nl�	�Пc[164[w��5�9[x�qG�y��tC8�|�29��o�%�1� ��{��m��!���� �0�B���f�x�����0����o���80��@'9K~���2P �����\�� '9K����@��������1��@/$/6/H/Z/U�|�?ainedi'ߑ/�/�/�/�/P�co�nfig=sin�gle&|�wintp���/$?6?H?Z?�	�ߐ??ٷ�gl[57�ٳq��?�;gp�08�ݲ07I�?F4��F2JO[6�:�?`)O�O�x �� �4s�x�O���$�� `�o�H_Z_l_~_�_�_ Q��_�_�_�_o o�_ DoVohozo�o�o�o�!�;�$doub5o���13��&duaml�i38��,4�o&�o9�o�n�o�a 8���Ao���P�&�8��%3L=}!��o�b8@������� ��z���(�:��+y:T��i48,2o�`�b{����ʟ {? �;�M�sc���;���As�� �}���e�u��X��@�F7L���`꠾O��2�h�z�6e�u7�����ｿϿ���̏�27��G�Y� k�}Ϗ��0�s����P�����!�1� M�_�q߃ߕ������ �������7�I�[� m����������� ���!�����6(�]��o��������$��74�6�����)�C��ߟT�	TPTX�[209�<Aw2 IHJ���Bw1H�@]H�����0�2��A#��[TtAv`��O�L#_�0�� \��5S[�treeOview3v�3��~~�381,26 M/_/q/0�/�/�/�/ �/�/~/?%?7?I?[? m?�o/(��o5%���?L�?�?�A�?\1~��?8"2��eOwO�?�? (}�LEK��O�O_�O ��8@�ONOa_s_�_��6_d�E_�_�_�_o V�#_���_�Sooo�o �oB�o�o��oA�o q+=Oas ��o������ �(�9���Q�x����� ����ҏ?����,� >�P�ߏt��������� Ο]�����(�:�L� ^�ퟂ�������ʯܯ k� ��$�6�H�Z�� l�������ƿؿ�y� � �2�D�V�h����� �ϰ������ϕo�o� �o@ߧE�c�u߇ߙ� �߽�����O����)� <�M�_�q���W��� ������&�8���\� n���������E����� ��"4��Xj| ����S�� 0B�fx�� ��O��//,/ >/P/�t/�/�/�/�/ �/]/�/??(?:?L? ��߂?1ߦ?���? �?�?�?O$O5OGO�? SO}O�O�O�O�O�O�O �O��2_D_V_h_z_�_ �_�/�_�_�_�_
oo �_@oRodovo�o�o)o �o�o�o�o*�o N`r���7� ����&��J�\� n���������E�ڏ� ���"�4�ÏX�j�|� ������a?s?蟗?� sO_/�A�S�e�w��� ������������ ,�=�O�a�#_������ ο��=��(�:�L� ^�pς�Ϧϸ����� �� ߏ�$�6�H�Z�l� ~�ߐߴ��������� ��2�D�V�h�z�� ����������
��� �@�R�d�v�����)� ��������ƚԔ�*defaul�t%��*level8�ٯw����? tpst�[1]�	�y�tpio[23���u���J\�menu7_l�.png_|1	3��5�{�y4�u6���// '/9/K/]/���/�/�/ �/�/�/j/�/?#?5?�G?Y?k?�"pri�m=|page,74,1p?�?�?�?��?�?�"�6class,13�?*O<O NO`OrOOB5xO�O �O�O�O�O�#L�O�0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]ooo�o�`�$UI_US�ERVIEW 1�֑֑R? 
���o��o�o[m�o'9 K] ����� l���#�5��oB� T�f������ŏ׏� ����1�C�U�g�
� ��������ӟ~���� �v�?�Q�c�u���*� ����ϯ�󯖯�)� ;�M�_�
��~���� ��ݿ���%�ȿI� [�m�ϑ�4ϵ����� ���Ϩ�
��.ߠ�i� {ߍߟ߱�T������� ��/���S�e�w�� ��Fߨ����>��� +�=�O���s������� ��^�����'�� ��FX��|��� ���#5GY �}����p� ��h1/C/U/g/y/ /�/�/�/�/�/�/�/ ?-???Q?c?/p?�? �??�?�?�?OO�? ;OMO_OqO�O&O�O�O �O�O�O�?�O_ _�O D_m__�_�_�_X_�_ �_�_o!o�_EoWoio {o�o0h