��   :�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����FSAC_LST�_T   8 �$CLNT_N�AME !$�IP_ADDRE�SSB $ACC�N _LVL  �$APPP  ����$8 AO  ����z�����o VERSI�ONw � 0��IRT�UALw�'DE�F\ � � �� ����ENABL�E� ������L�IST 1 �?  @!�,2��)����(y L^������ �-/ /Q/$/u/H/Z/ �/~/�/�/�/�/�/? �/:? ?q?D?V?h?�? �?�?�?�?O�?7O
O OmO@O�OdO�O�O�O �O�O_�O3___T_ <_z_`_�_�_�_�_�_ �_�W