��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� � P�COUPLE,  o $�!PPV1GCES C G1�!��PR0�2	 � $SOFT��T_IDBTOT_AL_EQ� Q1�]@NO`BU SPI�_INDE]uEX�BSCREEN_��4BSIG�0�O%KW@PK_F�I0	$TH{KY�GPANEhD� � DUMMYE1d�D�!U4 Q�*�0RG1R�
 � $TIT1d ��� 7Td7T� �7TP7T55V65V7*5V85V95W05W>W@�A7URWQ7UfW1pW1zW1�W1�W 6P~!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$^Nb_OPT�3�(�CELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1�UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t�d��MO� �sE 	� [M�s��2�wREV�BILF��1XI� %�R 7 � OD}`j��$NO`M@�+��b�x�/�"@u�� ����QX�@}Dd p E �RD_Eb��$�FSSB�&W`KBoD_SE2uAG� G�2 "_��B�� V�t:5`ׁQC ��a_EDu � �� C2��`S̐p�4%$l �t$�OP�@QB�qy�_�OK���0, P_C�� y��dh�U �`LACI�!�a���� �FqCOMM� �0$D��ϑ�@�pX��O�RB�IGALLOW� (KD2�2�@VAR5�d!�A�B e`BL[@S �C ,KJqM�H`S�p�Z@M_O]z��w�CFd X�0�GR@��M�N�FLI���;@UI�RE�84�"� SW�IT=$/0_No`S��"CFd0M�{ �#PEED��@!�%`���p3`J3t	V�&$E�..p`|L��ELBOF�  �m��m�p/0��C	P�� F�B����1x��r@1J1E_y_T>!Բ�`��gt���G� �0WARNMxp�d�%`�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�M�� R�r$OR�I�.&ӧRT�S�Fg CHGV0I��p�T��PA�I
{�T�P��� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8��9�4��x@�2� @� TRQ��$�%f��ր����_U���ѡ�Oc <� ����Ȩ3�2�ЯLLECM�-�MULTIV4�"$��A|
2q�CHILD>��
1��z@T_1b w 4� STY2�b4�=@�)24��8��@�� |9$��T�A�I`�E��e�TO���E��EX�T���ᗑ�B��2�2�0>��@ ��1b.'��}!�A�K�  �"K�/%�a��8R���?s  =�O�A!M��;A�֗�M�� 	�  =�I�" L�0[�� R�z�pA��$JOBB�x�����TRIGI�# dӀ����R��-'r��A�ҧ��_M���b$ tӀFL�6�BNG�A��TBA� ϑ�!��
/1�@À�0���R0�P/pX ����%�|���Bq@W�
2JW�_)RH�CZJZ�_*zJ?�D/5C�	��ӧ��@��Rd&A������ȯ�qGӨ�g@NHANC��$LG/��a2qӐ� ـ�@��A�p� ���aR���>$x��?#DB��?#RA�c?#AZ�t@�(.�����`FCT����_F࠳`�SM��!I�+lA�% ` �` ���$/�/�@���[�a��M�0�\��`��أHK��A�Es@͐�!�"W��Nz� SbXYZW�`�"����6	���I��'  �. II��2�(p�STD_C�t�1Q��WUSTڒU�)#�j0U[�%?IO1���� _Up�q�*c \��=�#AORzs 8Bp;�]��`O6  RSY�G�0�q^EUp���H`G�� ��]�DB�PXWORK�+~* $SKP_�p؂�A�TR�p , �=�`����Z �m�OD3��a _C`"�;b�C� �GPL:c�a�tőS�D�W�3Bb����P�.�� )DB�!�-,�B APR��
I�Ja3��. /�u���.����LuY/�_�����0�_����PC�1�_���r~�EG�]� 2�_��SVPRE.��R3�H $C��.$L8c/$uSނz �IkINE�WA_D1%�ROyp��������q�c7 t@�fPA����RETURN\�b�MMR"U��vI�CRg`EWM@^�SIGNZ�A ����e� 0$=P'�1$P� m�2p�p'tm�+pD�@ �'�bdNa)r>�GO_AW ���@ؑB1I�CS,d�(�CYI�4���`�1w�qu��t2�z2��vN�}��E}sD�EVIs` 5 oP $��RB���I�wPk��I_#BY���"�T7Q�t�HNDG�Q6 �H4��1�w��$DSBLC��o��vg@4��|tL��7O�f@�]���FB���FE�ra8�ׂ�t}s���8�> i�T1?���MC�S���fD �ւ[2H� W��EE���%F�p���t����9 T�p<��x�NK_N:���j��U��L�wHA�v	Z' ~�2���P~r��q7: �=MD	Ln��9�ጂٱh�����!e����J ��~�+����,�N�D����3��ՒG!aq�SLAd�7;  ��INP��"�����X}q_ �4<�06`�C� NU��  jD�Lק��SH!�
7=M��q���ܢ�Ӣ���g���>P +$ٰ�٢���^��^�Y�FI B\��Ă��'A	r'AWl�NTV��r]�V~�X�SKI�#�T���a�ۺ�T1J�3:3_�P�SAF�N���_SV�EOXCLU��N@�%DV@L��@�Y����S�HI_V
0\2P�PLYPRo�HI�M�T�n�_MLX�>�pVRFY_�ClM��IOC�UC!_� ����O�qţLS�0v�FT4Q������@P�E$t�t��A��CNFt��6եu��pm�4ACH�D�o������AF&C CPlV�TQTP8?�� �� ?`�@�TA�@�0L@ r��N��]� @����T��T! S����t<e@{RA DO�� �w2���!$n��_1�#�H!�̔��΀K��B�2��M/ARGI�$����A ��_SGNE�C;
$�`�a ^aR0��3��@ B��|B��ANNUN�P@?���uCN@�`�%0����� ���BEuFc@I�RD @Q�1F���4OT�`�s�FT�HR,Q��CQ0�M��NI|RE���r��AW���DAY=CLOAD�t;T|�<S�5}�EFF_AX�I��F`1QO3O���Eq��@_RT+RQE�G����0+RQ�2Evp ��|�F�0f�R0 ��tM�AMP�E><� H 0�``œ^�`Ds�DU�`����BCAr� �I?�`N ErID?LE_PWRI\4V!n0V�wV_[ |྅ �DIAG�5J�� 1$V�`SE�3TQl�e��0Pl�^E_��Y��VE� �0SW�H�q(� �b|�G�n�OHxPPLHZ�IRAl�B�@ �[��a�b�1�w3��O � ��v�|�I��0 �pRQDWf�MS-�%AX{<6Y�LIFE�@�&�MQy�NH!Q%��$F#C����CB0��mpN$�Y @�aFL�Al���OV0]&H�E��l�SUPPO$�@u�y��@_�$�冀!_X83�$gq�'Z�*W�*B1�'T�#`�fk2XZáY�Y2D8ECY`T@�`N����f� �C�I2���ICTA�K `�pCACH�ӫ�3з���I��bNӰUFFI� \��@���;T��<S6CQ.�MS�W�5L 8	�KE�YIMAG�cTM La��*Ax�&E���B��OCVIER-aM; ��BGL����y�?� 	��П4�N�:�ST�!�BP�D,P�D��D<��@EMAI䐔a���M�r�FAUL�|RObB�c�� spU�ʰMA"`T'`E�PO< $S�S[ v� ITw�BUF�7�y��7�tN[�LSU	B1T�Cx�o�R�tRSAV|U>R'c2 �\�WT���P�T�*`Sn�_1PbU���Y�OT�bK��P��M0��d���WAX��2�b��X1P��S_GH#�
��YN_���Q� <Q�D��0����M�� T�F��`|�\�DI��EGDT_Pɰ:�R��b�GRQM�&��Jq�a����׀��Fs� 7S (�SVqpB���4�_�.��a��T� �@���B�S7C_R]1IK>B'r��$t��R"A#u�H�a'DSP:FrP�lyIM|Sas�qz��a� �U>w� <1%sM�@I�P��s��0`tTH�b0ЃTr��T`asH9S�cCsBSCʴq0�� V�����S�_�D��CONVE�G ���b0^v1PFHy�adCs�`&a?ASC����sMERg��aF�BCMPg��`ETn[� UBFU� DU%P�D�:12��CDWy�p�P�CG�&[@NO6�:�V� �H�� ���P���C�����w��A��`���WH *�L Ơ�Cc�W����Y�� ���р�q�|��񨀖A��7}�8}�9P}�H ���1��1��U1��1��1ʚ1ךU1�1�2��2�����2��2��2��2�ʚ2ך2�2�3J��3��3����3��U3��3ʚ3ך3��3�4��QEXT[�X[b�H``t&``�z�k`˷$���FD�R�YTPV���RK"	��K"RE�M*F��]"OVM�:s/�A8�TROVf8�DT�PX�MXg��IN8ɉ W��IN	Dv�H2
�ȕ`K ^`�G1a�a��@Q%7Da�RIV��u"]"oGEAR:qIO.	K(�H4N�`���,(��F@� I3Z_MC�M<0K! �F� U�T���Z ,�TQ?' b�y@t�G?t�E |�.�>Q����[ �Pa� RI�E���UP2_ \ ��@=STD	p<TT����������a>RBACUb] T��>R�d�)�j%C�E��0��IFI��0��i�{�4��PTT��FLUI�D^ �?0gHPUR�gQ�"�r�a��4P+ I�$��S�d�?x��J�`C9O�P�SVRT��N�x$SHO* ��CASS��Qw%�pٴBG_%��3�����FORCx�B��o�DATA��-_�BFU_�1�bb�2�am=mm�b0��w` |��NAV	`�������$�S��Bu#$VISIl���2SC	dSE������V��O�$�&�BK�� ��$�PO��I���FMR2��a ��	��`# ��&�8�O� (��_����+IT_�^�ۄ)M�����D�GCLF�DGDMY�LD����5Y&H��Q$Y�M됇CbN@�{	 T�FS�P�Dc P��W�c>K $EX_WnBW1%`]��"X3��5��G+�d Y���SWeUO�DEBUG��-��GR��;@U�BK�U��O1R� _ PO_ )����:�M��LOOc>!SM� E�R�a��u _E e >@~�G�TERM`%}fi'�ORI�are gi%y�SM_�`�>Re hi%V�(i�i%3UP\Bj�3 -���e��w#�� f��G�*EL�TO�A�bF�FIG�2�a_���@�$�$�g$UFR�b�$�1R0օ� OT�_7F�TA�p q3N;ST�`PAT�q�0��2PTHJ�ԀEt�@�c3ART�P�'5�Q�B�aREL<�:�aSHFT�r�a�1�8_��R��у�&% � $�'@i�
�8���s@bSHI�0��Uy� �QAYLO �p�Oaq�����1����pERV��XA�� H��m7�`�2%�P�E�3�P�RC���AScYM�a��aWJ07����E�ӷ1�I��ׁUT�`Oa�5�F�5aP�su@J�7FOR�`�M  �O!k�]��5&�0L0��`H9OL ;l �s2T�,���OC1!E�$OP��qn�F��$�����$�2�PR^��aOU��3e��R�5e�X�1� �e$PWR��IMe�BR_�S�4��� �3�aUD��k�Q��dm��$H�e!^�`ADDR˶HR!�G�2�a�a�apRR\��[�n H��S�� ��%��e3��e���e��cSE��z�HS�;MNu�o���P0ªq��0OL�s߰�`ڵ�I ACROx��&1��ND_C�s���AfdK�ROUP���R_�В� �Q1 |�=�s���y%��y-���x���y���y>�=Ax��Ҁ�AVED�w�-��u&sp $���P_D�� ��^'rPRM_���!_HTTP_�H[�wq (ÀOBJ��l�b �$˶LE~3���\�r � (���ྰ_��TE#ԂqS�PIC��KRLPi?HITCOU�!��L���PԂ������PR��PSSB�{�J�QUERY_FL�Avs�@_WEBS;OC���HW�#1��s�`<PINCPU(���O���g������d��t��O� ��IOLN�t �8��R��$S�L!$INPU�T_U!$`��Pn G֐SL.�
��u���2�.��C���B�IOa�F_�AS=v�$L+ਇ+�A��bb41`�����Z@HYʷp����#qe�UOP:w `v�ϡ˶�¡�������"`PIC`����� �	�H�IP_sME��v�x Xv�cIP�`(�R�_N�p�d���Rʳp�ױ�QrSP �z�C��B�G(�� ��M�Av�y3 lv@CTApB��AL TI�3UfP_ l۵�0PSڶBU_ ID� 
�L � `�0Q0����0z)����ϴ�NN�_ O���IRCA_CN�f� { �Ɖ6-�CYpEA���� ����IC�ǫ�tpR<�=QDAY_
��NTVA�����!�8�5����SCAj@��#CL�
����
����v�|5�VĬ2b�l�N_�PCV�n�
���w�})�T��S�����
���e���T� 2|C Ր�� �v�~�8�֣�ذLAB1��\_ ��UNIX���� ITY裪��e~��p�� ��<)���R�_URL���$A;qEN ���s`vs�TeqT_U��m�iJ��X�M�$���E�ᒐR祪�� A��,���JH���FL�y��= 
���
�wUJR|U� ���AF�6G��K7��D>��$J7�s��J8B*�7���3�E�7���&�8\�)�APHI�Q4�y�DkJ�7J8R��L_K�E'�  �K�͐LMX� � �<U�XRi�����WATCH_VAZqxu@AំFIEL`�b�cyn���:� � bu1VbwPCTX�j�Y �LGE�߄� !��LG_SIZ΄�[8XZm�ZFDeIY p1!gXb ZW �S `�8�m��� ��b ��A�0_i0_�CMc3#�*'F Q1KW d(V(Bbpo pm�p� |Io�1 p�b pW RS��0 7 (C�LN�R��۠�DE6E�3����c�i���PL�#�DAU"%EA`q�͐�T8". GH�R���y�BOO�a��� C��F�IT0V�l$A0��RE���(GSCRX����D&�|ǒ�qMARGI� Sp�,����T�"�y�	S��x�W�$y�$���JGM7MNCHLt�y�FN��6K@7�r�>9UFL87@L8F�WDL8HL�9STPL:VL8"�L8s L8�RS�9HOPh;��C�9D�3R��}P�'IU h�`4�'�5$ ��S2G09�pPOWG�:�%`�3,64��N9EX��TUI>5I� �ӌ������C3�C<0'�@,�o:��&�@�!Naq�vcANAy��Q�A�I]�gt7Ӝ�DCS����cRS�cRROXXO"dWS�ÂRoXS{X�(IGNp 
Ђ=10 ܰ�[TDEV�7LLF��CZ!*�C �	 8�Tr$f/蛒h����3A�a�	 �W�萦�Oqs�S1Je2Je3Ja��BSPC � �ƋG`-T��%��Q�T�r@X�&E�fST�R9 �YBr�a �$E�fC�k�g��f	v8��CB� L���� � ��u�xs뀔�g�q��jt:�!�#_ ����ʐv�#Ӡ �s ��MC�� ����CLDP᠜�TRQLI ���y�t�FL���rQ��s5�D���w~�LD�u�t�u�ORG���1�RESERV��M����M�ŒC�s��� �� 	�u�5�t�uS�V��p��	1���>��RCLMC��M��_�ωА��: MDB�Gh�I����$DEBUGMAS��(����U�$T8P���EF�d�
�MF�RQҤ� � �K	HRS_RU��bq��A��$EFgREQUu!$0YOVER�k�t�f�PU1EFI�C%Gq�� �6�Y��z�� \����E�s$U�`��?���
�PSI`��	��C A ��ʲ�σUY�%��?( 	��MI;SC�� d��akRQ��	��TB� �� ���A��AX��𑧪�EXCE�Sg��d�M�H��9�u���9d�SC>�` � H�х�_�����������p�KE��+�� &�B�_, FLICBtB�� QUIRE CMEOt�O���r�LdpMD� �p{!��h5b����ND!���I����L �D|;
$INAUT�!�
$RSM�ȧPN��C�PSTL�H� 4U�LOCf�fRI"��eEX���ANG.R.���OD-A]��q��� �RMF0����icr�@mu���$�SUP�iu��FX��IGG>! � ���cs �F�cs
Fct��ޒ�b 5��`E��`T�5�tC�ьg�TI��7�Mܧ��� t��MD���)��XP��ԁ��qH��.���DIAa��Ӻ�W�!��0af���D@#)֡O�㥀�ෛ �CUp V 	���.����!_���� �{`�c������ |�P|��0� ��P{�KEB��e�-$B��o�=pND�2ւ����2_TXltXTRAXS���M���LO: ���L�}� ���C�.�&��RR2h��O� -�!A��� d$CALI����GFQj�2F`RsINbn�<$Rx��SW0ۄ���ABC��D_J��{�q��_J3��
��1#SP, �q�P�����3��H�9pq�#J��3n���O�QIM<�M�CSKP�zbH7?SbJ+�M�Qb��y����_AZ��/�EL�Q.ցOCMP��N�� cRTE�� �1�0 ����1��@ Z�SMG�0����J�G�pSCLʠ��SPH_�PM��f��zq�u�RTER��n�Pk�_EP�q²`A� �cM��DI��Q23UdDF�  ���LW�VEL�qINxr�@�_BLXP.��Y/��J��'$Q�IN���]�C�9%�".��8!6p_T� �@F%a"�6#a!��k)��Q�DHʠ��\�9`$Vw��_�A�$=����&A$���S�h��H? �$BEL� m���_ACCE� �	8�0IRC_4�q�@�NT��cO$PSʠ�rL���M4�s9 .7��GP@/6��9�7$3�73S2T�͡_Ga�"�0�1���8�1_MG}�DD�1���FW�p��3��5$32�8DEKPoPABN[7ROgEE�2KaBO�p�Ka���1�$US�E_v�SP��CTERTY4@� �� <qYNg�A�@�FR ��B�AM:�N�=R�0O�v1�DINC(��B��4���GY��ENC�L��.�K12��H0IN�bIS28U��O�NT�%NT231_���fSLO���|P��Iذ~��V�~� $��hpU#�CQ MVMOSI�1<�[�1���M�PERCH  �S��� �W���S lщR��l����E�0$�0PAS2EeL�DP�7�ONUЉZ�f�VT3RK�RqAY"�?c ��aS2�e�c�����BP�MOM�B��� C�H�}�Cj��c�3�gBT�DUX �2S_�BCKLSH_C S2Fu:��V���C-�es�Roz�A�CLAL�MJT@��`� �uCH�Ke ����GLRT�Ypн�8T��5���_��ùT_UM3��vC�3��1Z���LMT��_LG��%���0�E*�K�=�)�@5F�@8` 9�Nb��)hPC�Q�)hHТ��5�uCMqC���0�7CN_��1N���;SF�!iV�B��.W���S2/�nĈCAT�~SH�� ���4 V�q/q/V�T1���0PA�t�B_	P�u�c_f Z�f�P0e�cݔ�uJG����ѓ�OGއ�TORQU~@�S�i @`e��R� @B�_Wu �d�!a��#`��#`�UIh�Iv�I�#F��`S�:��I�0VC00��֢1ܮ�0���JRKܬ!���<�DBXMt�<�M��_DL�!_bGR�Vg�`��#`��#A�H�_%�?��0��COS��� ��LN#���ߥ Ŵ� ��=�������İ�<�Z���VA�MY�Ǳ:ȧ��᯻[�TH�ET0�UNK23��#���#ȰCB��C5B�#Cz�AS�ѯ�`�����#����SB�#���GTSkZAC�����&���$DU�phg6�j���E�%Q%a_��x�NEhs1K�t�� y�A}Ŧկ׍�����LPH����^U��Sߥ����������P!��(Ʀ�V��V��T� ��V��V��V
�UV�V&�V4�VB�H��������d�����UH
�H�H&�H4�UHB�O��O��Os����O��O��O
�O��O&�O4�O(�F��Ҫ�	���SP�BALANCE_lJ�6LE��H_}�SP>!۶^�^��PFULCb�q؉��K*1�UT�O_�p�uT1T2�	
22N�q2VP��M�a� i�Z23	qT�u`O�1Q�INSsEG2�QREV��PGQDIF�ep)1١U�1��`OBK�qj�w2,�VP�q~I�LCHWAR4B�"AB��u$MECH��J��A��vAX�aPo���׫"� � 
�?�10U7ROB�PCRS2#%�Ղ���C1_ɒT� � x $�WEIGH�@�`�$��\#��I�A�PI9FvA�0LAG�B��qS�B:�BBIL�%cOD�`�Ps"ST0s"P:�pt �!N�C!
L �P 
P2�Aɑ�  2��Tx&DEKBU�#L|0�"5�OMMY9C59N���$4�`$D|1 a�$0ېl� _��DO_:0AK!� <_ �&� �q�A���B�"� NJS�8_ԍP�@��"O�p _�� %�T7P�?Q�TL4F0TI�CK�#�T1N0%�3=p�0N�P� u3�PR\p�A��5��5U0_PROMP�CE��? $IR"��Ap�p8BX`wBMAIF�h�A�BQE_� OC�X�a�@RU�COD��#FU�@�&ID_��P�E82B> G_SwUFF�� �#4�AXA�2DO�7/�5� �6GR�#��D C�D��E��E-��D�U4� �_ H_F�I�!9GSORDf�! R 236s��HR�AN0$ZDT�E�P�!X5�4 =*WL_NA�1�0|�R�5DEF_I�X �RF�T�5�"�6�$�60�S�5�UFISm�#� m1|��40c�3�T6�"44􁆂�"D� ?r�fd�#D�O@ l2LOCKE���C�?O0G2a�B�@UM�E�R �D�S�D�U�D>b�B�c �E�S�Dd�B�&2v2a �C�ʑ�E�R�E�S�C9wwu�H�0P} d�0�,a��F0W�h�u�cΐ �TE�qY4�� �!LOMB�_�r�w0s"VIS���ITYs"AۑO>�#A_FRI��F~SI,a�n�R�0H7��07�3�#s"W�!W�Q��%�_���AEAS{#�B��|��x`WB8�45�55�6�|#ORMULA_�I���G�W� �h 
>75COEFF_O�1&)�$�1��Go�{#S� 52�CA� :?L3�!GR�m� � � �$�`�v2X�0TM��g���e�2�c��3E�RIT�d�TAP� M �LL�Dp`S��g_SVkd��$�v�AP�.���AP� ޅ�SETU,cMEAG@�@Πt �!HRL �� � (�  0��l��l��aw�"�R�0�a�a}d]�Ad��B��Ay`Ga�x`��[Ѐk@RE�C[Qq��1SK_�A y�� P_!1_USER���p�*���VEL�� ��-�!��IzP� w�MT�1CFG����  �0]O�NOREJ �0l����[�� 4 �e���"�XYZ�<S�� 3� ��_7ERRK!� U ѐ�1�@c�Ȱ�!�>��B0BUFINDqX���p� MORy�7� H_ CUȱ�1���dAyQ?�I>Q'$ +�a������ \�G{�� � $SI�h��@�2	�VOv�q�- O�BJE| w�ADJ1UF2yĈ�AY�����D��OUKP���\�AMR=�Tp��-���X2DIR�����Xf�1  DYNHt�0�-�T� ��R���0� ���OPWO}R�� �,B0�SYSBU����SCOPo���z�Uy�bXP�`K���PA��q������OP�@U����}�"1��IMAG۱_ �п"3IM.���IN����~��RGOVRD"���	���P����  >PgplcC��L�`BŰ|?l�PMC_E�P�1N��Mr�12112R�"�SL| ���� �R OVSL:=S�rDEX\a`"��2�:�_"��� P#���P������2�C �P>���#�/_ZERl���:����� @��:��O&�@RIy��
[�g@�e���s�P�PL����  $FREEY�EU�~�Z���L����T�� A�TUSk�,1C_T�����B������p��Vc1��P��� Dc1�к���LQ����0MQ��ۡL�XE��x�5IP�W�` ��cUP��H`&aPX;@���43�� ��PGY��g�$S�UB���q���J?MPWAIT~ ���LOW���1wē �CVF_A�0��RX�Z��CC �R$���28IGNR_P�L��DBTB� P�*a�BW@.t�UL�0-IG��!@I�OTNLN,�RB��b�N!@��PEE�D~ ��HADOW� ��t���E�����ܹ�PSPD��� L_ A�нP���	#CUNq � �RP F(�LYwPa����_PH_PK���b�?RETRIE��x������� H�0NFI���� ���V �$ �2�d�DBGL�V<LOGSIZ,z�baKTU���$�D��_TXV�E�M�Cڡ��� �-R��#�r��CHECK�z����L���ϰ�q)�L��NPAB�`TJ"����)1P����
�AR�"�BC �=Sa��O�@����ATTS�u䡳&� w�^a�3-#UX^�4�sPL�@Z�� $d�~�qSWITCH�Zh�W��AS��f��3LLB���_ $BA�Dvc��BAMi��6I��(@J5��N�UB6|[F
A_KNOWK34qB"�U��AD+Hc�� D��IPAYL#OAq�9p�C_���GTrѼGZ�CLqAj���PLCL_6� !4��BOA?�T7�VFYCӐ�Jp��D�I�HRՐ�G粒TB��6�J��zQ_�J�A �B�AND�����T�BQ�q��P�L@AL_ �@�0 =�TAe��pC��uD�CE���J3�P��V� T�PDC�K^�)b��COM�_�ALPH�ScBE0<�߁�_�\�X�x>\� � ���OWD_1�J2�DDM�AR<�h�e�f�cQѯTIA4�i5�i6��MOM(��c�c�ch�c�cV�B� AD�cpv�cv�cPUBP�R�d<u�c<u�b}"�1����� L$PI$��pc��G�y�T�I�yI�{I�{I�s��`�A���v��v��J�b��a��HIG�3���0��� 5�0�f�?�5N�5�SAMPD Ƣ��0����;@�S  ��с6���1���� � ��`���`1�K�P��`�腽P�H��IN 1��P��8�T�/��:��z�Q�z���GAMM�&�S��$GE�T�����D^d>�
�$�PIBR��I.��$HI��_���$1��E=��A�9�*�LW�W�N�9�{��*�Zb���QCdC�HK0�j�ݠnI_��M�JļRoh�Q ���sJ�-v��S ��$�X 1��N�I�RCH_D$RN���^�LE��i�p�Zh8�}ţMSWFL/�M�PSCR�75�Ҽ ��3�"Ķ�6���`��ع�紙��0SV��P'�������GRO�g�S_�SA=AH�=ńNO^`Ci�_d=��no �O�O�x�ʚ��p�B�u,�ȐcDO�A��! �ں�*�t�:�Z1f��;�7����C etM�mu� � �YL�snQ ��� ���"��<s�	������nQ૰<3M_Wl�����\p��(�oсMC��P���Q ����hpM.�pr�� ��!��$�W<M��ANGL�!�A M�6dK�=dK�DdK��TT7�Nk@��3�#�P%XC OEc�QZ��hp�	nt� ���OM���ϑϣϵ���p�`� c�Z0���hp:^a_�2� |a� J��i���c���cJ��j �����jA�{ �{�J��{ �@{�P�1��PMON_QU��� � 860Q�COU��QTH�xHO��B HYSf�0ESPBB UE- t3�f0O�4�  c �P�^�RUN_+TO��gpO���� P�@��I�NDE�#_PGRA����0��2��NE_3NO��ITf��^o INFO��a"h�����H�OI�� (*�SLEQ�!�*�*�Q OS���l4� 460E�NABy� PTION�3��r��^wGCF�!� @60�J�Q���R��d!��u�PED;IT�� �� ��KAQ"� �E(�N9U'(AUTY�%COPYAQ�2,�q�e�M�N< @+��PWRUTm� C"N�;OU�2$G��$�
�RGADJ��u2X_��IX����&���&W�(P�(~��&�9�� 
�N�P_CY�Cy�w�RGN�Sc�{�s�LGO�£�NYQ_FREQSrW@��X1�4�L�@�2P0�!�c@��"�CRE��MàI�F�q�NA��%��4_Gf�STAT�U~�f��MAIL䩂|CIq�=LAS�T�1a*4ELEM�g� ��QrFEASIt;�ւΰ���B"�F�AF����I � ��O2�E u�vB�AB��PE� =�V@A�FzQ�I��TqU[���R��S�FRMS_TRpC�Qc��C`��Z�
��1�D � �,2ns؆�	MB 2� `���N� 3V�R2WR*���шR8^W�wj�DOU�^��N�,2PR`�hٞ1GRID��B7ARS!�TYuB�OTOp�� �|_�4!� �R�TO|��d� � ����POR�c~vb�SRV�0)"dfDI[�T�`;aNd�pXgD
�Xg4Vi��Xg6Vi%7Vi8:a�Fʒg��z $VALU��C0�3D1@(1F05�� !pf���S1�1-ȆAN/��b��1R�]11ATOTcAL����=sPWE3�I�QStREGENQzfr��X�H�]5	�v( TR�CS�Qq_!S3��wfp�V�!��r��BE�3�PG0B��( sV_H�PDqA(��p�S_Ya����i6S��AR(�2�� �"IG_S!E�3�pb�5_� �t{C_�V$CMPl��DEp�G���IBšZ~�X�
�% Fm��HANC.� �p Qr�2���I#NT9`cq�F����MASK�3�@OVRMP �PD�1-�D�W� ��aХT�l�_RF�{�V�PSL)GP�g�9�j5��,�;pDpS���4���U���|�TE���`���`k����J^�Y�y3IL_M`x4�s��p��TQ( ����@����V.�CF<�P_ �R�F�M]�[V1\�V1j�2y�U2j�3y�3j�4y�4j���p۲�������ܲIN�VIB�8�6�#��*�2&�2�2�3&�32�4&�4�2��6�|�J�  ��T $MC_F,K `� �L>�J�х1pMj�Iу��zS� ��1���KE�EP_HNADD"��!鴓@�C��0A	��Q����
�O!��v ���p
�և
�REM!�	�Cq�RF��]�b�U�4e	�HP�WD  �S�BM���PCOLL�AB*�p��/q�2�IT/0��""NO1�FCALp⎵��7� , �FLv�A�$SYN���M���Ck��RpUP_�DLY��zDE�LA9�Dq�2Y A�D(��(0QSK;IPO�� �`� �O��NT����c�P_� ��׾ ��cp�� �q�����o`��|`�� �`�ږ`�ڣ`�ڰ`��=9�!�J2R0  �lX�@TR3H�� 1AH� �H���$ �RDCq��� �� R�R, 5��R��1��E��5TRGEp�_C��RFLG"����W�5TSPC��1UM_H��2/TH2N}Q�;� 1� y�E�D�Q02 � D� ˈ��@2_PC�3W�S���1Y0L1w0_Cw2$C+�n�� � $\�  U@��V7����� 0��� c�\���� � rd��C�Q,��7��DZ Gs�RUV�L1[�1h���10]�_DS�������PK 11�� l�ڰ����q��AT ?��$�Q[7�� ���K 5T���HOMME� *�c2h�n�����]�
`3h���!\3E `4h�hz�����5h���	//-/?/W6h�b/t/�/��/�/�/ ���!7h��/�/??'?9?
�8h�\?n?�?�?,�?�? _S����  �Aa{p���3�+�_�Ed�� T=�nD4vnCIO�䑎II@`�O��_�OP�E�C.rfBXP�OWE	�� �X@�f��$�$Cd�S�����_���3�3� ��@�SI��G�P0�QIR�TUAL�O
QAA�VM_WRK 2� 7U �0  �5�Qn_zXk_�] �\	�P�]�_3�8P!��_�_�Ve�\#m�/o�Q5ojo|o�dHPB�S�� 1Y�? <Xo�o �o�o�o#5GY k}������ ���1�C�U�g�y� ��������ӏ���	� �-�?�Q�c�u����� ����ϟ����)� ;�M�_�q����������˯ݯ�bC$�AXL�M�@iAQ��c  �d�IN����P+RE
�E�J�-�'_UP��[�7QHP?IOCNV_��k �	�Pr�US>��g�cIO)�V 1]U[P $E`��Q0ս9lҿ8P?��i@ ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o�o�o�o�m�LAR�MRECOV �a��-���LMD/G ��ɰ��LM_IF  ���ை����z�v���%�6�, 
 6�_��r� ��������̍$w��� ׏��8�J�\�n�����NGTOL  �a� 	 A �  ��ț�PPI�NFO ={� <v����1��  I�3�a�"rP��� t��������ί���>�o����j�|��� ����Ŀֿ������0�B�PzPPLIC�ATION ?����J��HandlingTool ��� 
V9.30�P/04ǐM�
�88340�å�F90����202�ť�|�Ϭ�7DF3���M̎�NoneM��FRAM� �6��Z�_ACTI�VE�b  sï� � p�UTOMO�Dz�A���m�CH�GAPONL�� ���OUPLEDw 1ey� �������g�CURE�Q 1	e{  T*���	p��xw���#r�g���e�HN����{�HTTHK)Y��$r��\[�m� ���O�	�'�-�?�Q� c�u����������� ��#);M_q ������ %7I[m� ��/���/!/ 3/E/W/i/{/�/�/�/ ?�/�/�/??/?A? S?e?w?�?�?�?O�? �?�?OO+O=OOOaO sO�O�O�O_�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q��c���1�TO��|��p�DO_CLEA�N��n��NM  �� �B�T��f�x���%�DSPDgRYR��m�HI���@/�����,�>� P�b�t���������ίj�MAXa�ۄ�������Xۄ������p�PLUGG��܇�Ӯ��PRC��B�" ��ׯF�OK���^ȔSEGF��K�� �����.�����,�8>�v���LAPӟ� ��Ϥ϶��������π�"�4�F�X�j߯�T�OTAL�7���U�SENUӰ�� ����ߖ�1�RGDI_SPMMC����C����@@Ȓ��O�ѐ�����_STRING 1
�ۿ
�M��S�l�
A�_ITE;M1K�  nl�g� y������������ 	��-�?�Q�c�u����������I/O SIGNALE��Tryout� ModeL�I�np��Simul�atedP�Ou�tOVER�RА = 100�O�In cyc�lP�Prog� AborP�~��StatusN��	Heartbe�atJ�MH F�aul��Aler�	�������*<N`  ׃G�ׁY�c��� ��////A/S/e/ w/�/�/�/�/�/�/�/wWOR��G�-1� ?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO�cOuO�O�O�NPO E��@E;�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8oJo�BDEV�Nu`�O bo�o�o�o�o�o�o ,>Pbt�������PALT��E?�A�S� e�w���������я� ����+�=�O�a�s����GRI�G뽑 1������	��-�?� Q�c�u���������ϯ�����)�����R �a�՟;��������� ѿ�����+�=�O� a�sυϗϩϻ���O�PREG��y��� -�?�Q�c�u߇ߙ߫� ����������)�;��M�_�q����$AR�G_-0D ?	��������  	$���	[��]���������SBN_CONFIG���� ��CII�_SAVE  ���)���TCEL�LSETUP ���%  OME�_IO����%M�OV_Hn�����R�EPd�����UTO/BACKY���#�FRA:\��� ����)�'`rl ��&� 7�"� 24�/06{  09:_35:24������͓����� �+=Oas��������� �/1/C/U/g/y/�/ /�/�/�/�/�/	?�/ -???Q?c?u?�?�?p�ׁ  _��_\�ATBCKCTL.TM���?�?�?O\ O��INI�Y��-���MESSA�G9�GA)��RKODGE_Ds�<��zH�Ow`�O��PAUS��@ !��� , 	�����O�G,		�O__ ?_)_;_u___�_�_�_ �_�_�_�_�_)m�D�@?TSK  �M&<,O��UPDT�@EG�d�`�FXWZD�_ENBED��fS�TADE��e��XI�S�UNT 2t��&�(�� 	\`��h� Q�� ��Q`)�3�����ʮq  Cp�Y,t:
p�5p�JUg~q�|P t����E3�����D�m�w%�G����aM�ETc�2LfE� �P qBb�B��B�B5RB��GB���CM�\��}?yo�?�٥@?��=@�u�?z�R@�i���}SCRD�CFG 1��� �A�&� �����ԏ�����Q=���H�Z�l�~� ����	�Ɵ-������ �2�D���域���G�R�`�`�O���0NA�����	��_�EDC@1n�� �
 �%-�0EDT-q����%�p��òu���������������  ����2����*�R�bB���*�q��������3bϮ�@Ͻϯd ?�����=�O���sϏ�4.ߞ�{�����W��� 	�߱�?ߏ�5��j� G����#������}�6��6��Z��΀��Z����I��7 �����&��λ�&m������8^ҿ����	͇�9K��o��9*�w�� 	�S��;��CR����B/T//��/��w//��РN�O_DEL����GE_UNUSE����IGALLOW� 1��   �(*SYST�EM*is	$S?ERV_GR�;B0n�@REGK5$m3i|B0NUMp:�3�=�PMU� iu�LAY�pi|�PMPALD@�5COYC10�.�>�0<�>CULSU�?�=��2�AM3LOWDB�OXORIt5CU�R_D@�=PMC�NV�6D@10|�>�@T4DLI�`�=O_9	*PROG�RAJ4PG_cMI�>�OPAL�E�_UPB7_B>�$FLUI_RE�SU�7p_z?�_�TMRY>h0�,�/�b�_ �_o o2oDoVohozo �o�o�o�o�o�o�o
 .@Rdv����������"L�AL_OUT �1;l���WD_A�BOR�0?d�IT�R_RTN  ����g�NONS�TOǠ�� 8CE_RIA_I0���ۀ��ŀF?CFG ��۔���_LIMY22�ګ �  G� 	i�J��<e�tg��5�� 9��������
���u���PAQPGP 1�����Q��c�u�4�CK0����C�1��9��@���PCV��CV��]��d���l��s��P���CU[٤m��v����}����� C�����-���?�ÂH=E� ONFI�Pq�nG�G_P�@1� �%��������ǿٿ����G�KP7AUSaA1�ۃ �2�W��Eσ� iϓϹϟ�������� ��#�I�/�m��eߣ���M��NFO 1�"��� ��7��ߖ��B���ƓA�&����ߌ��I��@�8� A�  %Cj��D����3���7�lB� 3�4E�ŀO��c�COLLECT�_�"�[�����E�N�@��y���k�ND-E��"�3�"�1234567890��\1�� �$�֕H&��)M�r� \,L�^���]+������ ������C 2� Vhz���� ��
c.@R��v�������΢� ����IOG !���q���`u/�/�/�/C'TR�K2"'-(׀^)
��.R�#R-�*W� 9�_MOR�$� �;�l5��l9�?r?�?@�?�?�;E2��%S=%,W�?@�@��C׀�K)DցC�R�&�u�XOWAWBC4  �A�q��׀x׀}A"@Cz  B�@�CG�B8��AC [ @yB�׀ց�:d�43 <#�
�E���I�O�C*=AI��'GM?�C��(S=���Qd=AT_�DEFPROG ��;%�/m_APINUSE�V�ۅ�T�KEY_TBL � s�ہ���	
��� !"#�$%&'()*+�,-./�:;<=>?@ABCDP�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������Ga�������������������������������������������������������������$��PL�CK�\���P�PST�An��T_AUTO�_DO��NFsI�ND���n��R_T1wT2N�����5ŀTRLCPLE�TE���z_SCREEN ��kcscÂU���MMENU 1)O� <�[_#� q��,�a���>�d��� t���ӏ����	���� �Q�(�:���^�p��� ����̟�ܟ�;�� $�q�H�Z��������� �Ưد%����4�m� D�V���z���ٿ��¿ �!���
�W�.�@ύ� d�vϜ��ϬϾ���� ��A��*�P߉�`�r� �ߖߨ��������=� �&�s�J�\����������'�,�p_?MANUAL�Eq�DB
12�v�iDB�G_ERRLIP9*�{h! 0��������g�NUML�IM�s:QOE�@D�BPXWORK 1+�{��>Pb�t��-DBTB_��q ,��kC3!�VD!DB_AW�AYo�h!GCP� OB=��A�_A!L���o�k�Y�p�utO@`�_�� 1-�+@
-k-6[�6�_M+pIS�`��@"@�ONTIM6�w�OD��&�
�U;MOTNE�ND�_:RECO�RD 13�{ y��[CG�O�f! T/[K��/�/�/�/_( �/�/f/?�/??Q?c? �/?�??�?,?�?�? OO�?;O�?_O�?�O �O�O�O(O�OLO_pO %_7_I_[_�O_�O�_ _�_�_�_�_l_!o�_ ,o�_io{o�o�oo�o 2o�oVo/A�o eP^�
��� R���=��a�s� �������*�ߏN�� �'���ԏ]�̏���� ����ɟ۟v���n�#����G�Y�k�}���TOLERENC�sB�0� L��g��CSS_CNST_CY 24	�t�	��.������ 0�>�P�b�x������� ��ο����(�:��äDEVICE ;25ӫ ��� �ϱ������������/�AߟģHNDG�D 6ӫ� Cz�T�.!ơLS 27t�S������������/�U�ŢPARAM 8Gb�A���Ք�RBT 2:.8�<����CkA� �~��  � A�p��.SB���~A�B�  ����������.`��  ����A�A�C����c�u����C�A�D��k�epz�A�A��HA�c��A�	�?(u�L^p���A�B�t/�D��C���_ 	 A=���ABffA#�33AҊ��ͳA�A�Cf��aĒ�A�J��7B]���B��B�ffBᴠ�33�C$.@R� ( ����A���� 
/��//)/;/�/ _/q/�/�/�/�/�/�/ �/<??%?r?I?[?m? ?�?�?�?�?�?&O8O �PObOMO�OqO�O�O �O�O�O_�OOL_ #_5_�_Y_k_�_�_�_ �_ o�_�_6ooolo CoUogo�o�o�o�o�o �o �o	h�O� w�����
�� .�	__I'�1_�q� �������ˏݏ�� �%�r�I�[������ ����ǟٟ&����\� 3�E�W����ȯ��� ׯ�"��F�1�j�E� s�����m�������ѿ �0���f�=�O�a� sυϗ��ϻ������ ��'�9�Kߘ�o߁� ����[����(��L� 7�p��m����� ������$�����l� C�U���y��������� �� ��	V-?� cu����
�� @+dO�s� �������*// /`/7/I/[/m//�/ �/�/�/?�/�/?!? 3?E?�?i?{?�?�?�? �?�?�?�?FO�jOUO gO�O�O�O�O�O�O_ _�'O9OO=_O_�_ s_�_�_�_�_�_�_�_ oPo'o9o�o]ooo�o �o�o�o�o�o: #5��O������ ��$��H�Fz��$DCSS_SL�AVE ;����w��~`�_4D  w����AR_MENU <w� >�؏� ��� �2�^rǏ\��n�\���SHOW �2=w� �  fr[q����Ə������,�>�D�b�t���  ����ҟϯ���� )�P�M�_�q������� ��˿ݿ���:�7� I�[ς�|Ϧ��ϵ��� ������$�!�3�E�l� fߐύߟ߱������� ���/�V�P�z�w� ������������ �@�:�d�a�s����� ������\���*�H� N�K]o���� ����28�G Yk}����� �"�1/C/U/g/ y/�/��/�/�/��/ /?-???Q?c?u?�/ �?�?�?�/�??OO )O;OMO_O�?�O�O�O �?�O�?�O__%_7_ I_pOm__�_�O�_�O �_�_�_o!o3oZ_Wo io{o�_�o�_�o�o�o �oDo-Se�o ��o�������.�=�O���CFG7 >�����q���dMC:\���L%04d.C�SV\��pc��������A ՃCH݀z@�v�w�#��q����:�J�8�7���GJP�j�)�́�p�+�n�RC_OUoT ?z������a�_C_FS�I ?�� |����� @�;�M�_��������� Я˯ݯ���%�7� `�[�m��������ǿ �����8�3�E�W� ��{ύϟ��������� ���/�X�S�e�w� �ߛ߭߿�������� 0�+�=�O�x�s��� ����������'� P�K�]�o��������� ��������(#5G pk}�����  �HCUg ��������  //-/?/h/c/u/�/ �/�/�/�/�/�/?? @?;?M?_?�?�?�?�? �?�?�?�?OO%O7O `O[OmOO�O�O�O�O �O�O�O_8_3_E_W_ �_{_�_�_�_�_�_�_ ooo/oXoSoeowo �o�o�o�o�o�o�o 0+=Oxs�� �������'� P�K�]�o��������� ��ۏ���(�#�5�G� p�k�}�������şן  �����H�C�U�g� ��������دӯ���  ��-�?�h�c�u��� ������Ͽ����� @�;�M�_ψσϕϧ� ����������%�7� `�[�m�ߨߣߵ��� �������8�3�E�W� ��{����������� ���/�X�S�e�w� �������������� 0+=Oxs�� ����' PK]o���� ����(/#/5/G/ p/k/}/�/�/�/�/�/� ?�/??H?C?U3��$DCS_C_F�SO ?�����1 P [?U?�?�?�? �?�?O
OO.OWORO dOvO�O�O�O�O�O�O �O_/_*_<_N_w_r_ �_�_�_�_�_�_oo o&oOoJo\ono�o�o �o�o�o�o�o�o'" 4Foj|��� ������G�B� T�f���������׏ҏ �����,�>�g�b� t���������Ο��� ��?�:�L�^����������ϯʯܯg?C_RPI~>�?�;� d�_�
�}?.�p����,ݿj>SL�@��� 9�b�]�oρϪϥϷ� ���������:�5�G� Y߂�}ߏߡ������� �����1�Z�U�g� y������������ 	�2�-�?�Q�z�u��� ����������
 )RM_q��� ����*%7 Irm���� �/�ϛ�,�/W/ �/{/�/�/�/�/�/�/ ???/?X?S?e?w? �?�?�?�?�?�?�?O 0O+O=OOOxOsO�O�O �O�O�O�O___'_ P_K_]_o_�_�_�_�_ �_�_�_�_(o#o5oGo poko}o�o�o�o�o�o  �oHCUg ��������� ����NOCOD�E @������PRE_C�HK B��3�A� 3��<� �7��������� 	 <�����?#ۏ %�7��[�m�G�Y��� ����ٟ�ş�!��� �W�i�C�����y�ï կˏ������A�S� -�_���c�u���ѿ�� �����=��)�s� ��_ϩϻϕ������ ��'�9���E�o�I�[� �߷ߑ���������#� ���Y�k�E���{� �����������C� U��=�����w����� ����	����?Q+ u�a����� �);_qg� Y��S���� %/�/[/m/G/�/�/ }/�/�/�/�/?!?�/ E?W?1?c?�?���? �?o?�?O�?�?AOSO -OwO�OcO�O�O�O�O �O_�O+_=__I_s_ M___�_�_�_�_�_�? �_'o9oo]oooIo�o �oo�o�o�o�o# �oGY3E��{ �����o�C� U��y���e������� ����	��-�?��K� u�O�a��������� ͟��)��1�_�q�� }�������ݯ�ɯ� %���1�[�5�G����� }�ǿٿ������� E�W�1�{ύ�G�u��� �ϯ������/�A�� -�w߉�c߭߿ߙ��� ������+�=��a�s� M���ϑ������ �'��3�]�7�I��� ������������� ��GY3}�i� �������C /y�e��� ����-/?//c/ u/O/�/�/�/�/�/�/ �/?)?�?_?q?K? �?�?�?�?�?�?�?O %O�?IO[O5OO�OkO }O�O�O�O�O_�O3_ E_;?-_{_�_'_�_�_ �_�_�_�_�_/oAoo eowoQo�o�o�o�o�o �o�o+7aW_ i_��C���� �'��K�]�7�i��� m��ɏۏ������ �G�!�3�}���i��� ş������1�C� �g�y�S�e������� ���ѯ�-���c� u�O�������Ͽ�ן ɿ�)�ÿM�_�9�k� ��oρ����Ϸ��� ���I�#�5�ߑ�k� ���ߡ�������3� E���Q�{�U�g���� ���������/�	�� e�w�Q����������� ����+Oa� I������ �K]7�� m�����/� 5/G/!/k/}/se/�/ �/_/�/�/�/?1?? ?g?y?S?�?�?�?�? �?�?�?O-OOQOcO =OoO�O�/�/�O�O{O �O_�O_M___9_�_ �_o_�_�_�_�_oo �_7oIo#oUooYoko �o�o�o�o�o�O�o3 Ei{U��� �����/�	�S� e�?�Q�������я� �����O�a��� ����q���͟����� ��9�K�%�W���[� m���ɯ�����ٯ� 5�+�=�k�}������ �������տ�1�� =�g�A�Sϝϯω��� �Ͽ�������Q�c�����$DCS_�SGN CS�����#M��01-AUG-2�4 15:42 |EӘ�6-JUN�џ09:39������� X�L�������������Д���M��Þ�ǧj�����{�VE�RSION ���V4.2.�10�EFLOG�IC 1DS���  	�D���X�k�X�z�M�P�ROG_ENB � ��b��Л�U?LSE  ����M�_ACCLI�M��������WRSTJNT�����w�EMO���ѷ�L��INIOT EZ�O���OPT_SL ?�	S�1�
 	�R575�Ӆ�74*��6��7��5A��1��2��l���G�h�TO  t���.�H�V?�DEX��d����FPATHw A��A\4����HCP_CLNTID ?+�b� l������IAG_GRP� 2JS�� �a[��D�  D�� �D  B�  ;B�@ff��/CB�@[��W�@��q��B�N��C�-Bz�w�Bp@e`���mp3m7 �78901234�56�*�[�� � Ao�mAj�1AdA]��
AW|�AP��AJ-AC�/A;�A4�H���@�  Aʩ�A�A3!_A�@@��B4��� ��t���
�u�ƨApffAj��yAeK�A_��AY��AS�� MC�AF��A@ �O�+/=/O$�O�c K�w(@�X�?8��@��y�/�/�/�/�/8��;d�2�5?@~�ff@x1'@q���@kC�@d��D@]��@Vv�6?H?Z?l?~?8�s�0l��@e���@^��@W\)@O��@H�0�?<@7K�@.V��?�?�?�?
O8S�@M00G<@A���@<1@5���@/l�@(�Ĝ@!�0�\ NO`OrO�O�Ox'g�L_ K�;_�_�__g_�_�_ �_�_o�_�_�_Yoko@Io�o�o+o�oX�"�� 2�17A�@J>���R
q?�33?wY��r��J�7'Ŭ2q63p4w�F>r��LJ�@�p�Zr�
=�@�@�Q�jq��@G Ah�@���@�T= c<���]>*�H>�V>�3�>����J<���C<�p�q�x��� ��?� �C� � <(�U�� 4Vr�33��@
���A@��?R�oD� �mR�x���Q��t�����Z�Џ��؏�,��i?��7N�>�(�y>�@Z�=���Jo��G�v�G�J �B�E�����a��@ǐ�@���@��@OQ�?L ���ŲI�P���&�
��'��@�K�����Ag�q�PC�  ?C���Cuy�
���ʯ ?����	��Ԡ��4���X��v����*A DCj��ZD C3���5�2B���F�ǿB��ֿ�����E�t�.�����x= �W�����P����S�3ϔ�	CT�_CONFIG �K3����eg��STB_F_TTS��
����"�������{�M�AU���MSW�_CF��L  �K �OCVIEWf	�MI�U��� �߭߿��������� �0�B�T�f�x��� ������������,� >�P�b�t�������� ��������(:L ^p����� � �6HZl ~������,/��RCB�N��!��F/{/j/�/�/��/�/�/��SBL_�FAULT O�9*^�1GPMSK���7��TDIAG� P��U�����qUD1:� 6789012345q2�q���%P�ϭ?�?�?�?�?O O+O=OOOaOsO�O�O��O�O�O �a6�I'�
��?_��TRECPJ?\:
j4\_�7_[�? �_�_�_�_�_�_oo (o:oLo^opo�o�o�o��o�O�O_ _�UM�P_OPTION��>qTRB���9�;uPME��.Y�_TEMP  ?È�3B����ps�A�pytUNI'���ŏq6�YN_BR�K Qt�_�EDITOR q&qh�r�_2PENT 1R�9)  ,&�MAIN �pNO� 0 TEIRA� &p5� &
P�EGA_%�b�&�PICK1_P�LACEW�8�&�L�BARRA_�ES��8�&C�OLOCA_bpA?_IRVIS$r�� &ЄPRE�NSA ޏ8�&SEGU������P�p�  &�-BCKEDT-� ��Q���C�PR�OG_1 [�m�SUMIR����>��DROP_DEsFE�p��ERT�����֜2�̟ޔ3��@�ЄANTEONA_C?�A�ؒ�SEMܕ �C��Є����Ƀx�UP��M4�<�������5�(��V���F+�D� ��F��E�T����%E�MGDI_STA�u~��q�uNC_I?NFO 1SI��b�������Կ�쮳��1TI� �P�o#��0�
0�d�o }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߯���������Hu�  �2�D�R�j�R�x�� ������������� ,�>�P�b�t������� ������Z��#5 Ga�k}���� ���1CU gy������ ��	//-/?/Yc/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?��?O%O 7OQ/GOmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �?Ooo/o�_[Oeo wo�o�o�o�o�o�o�o +=Oas� �����_�_�� '�9�So]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�K�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�C�5�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ��������!�;�M� W�i�{�������� ������/�A�S�e� w��������������� +E�Oas� ������ '9K]o��� �1����/#/= G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?��? �?	OO5/?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�?�_�_oo-O #oIo[omoo�o�o�o �o�o�o�o!3E Wi{����_�_ ����7oA�S�e� w���������я��� ��+�=�O�a�s��� ������ߟ��� /�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������͟ ׿����'�1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߫�ſ������� ��;�M�_�q��� �����������%� 7�I�[�m�������� ���������)�3E Wi{����� ��/ASe w��������� /!+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?/ ��?�?�?�?/#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�?�_�_�_ �_Oo-o?oQocouo �o�o�o�o�o�o�o );M_q�� �_����	o�%� 7�I�[�m�������� Ǐُ����!�3�E� W�i�{�����ß՟ 矝���/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߩ����� �������1�C�U� g�y���������� ��	��-�?�Q�c�u� ���߫����������� );M_q�� �����% 7I[m���� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?���?�?�?�?� OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�?�?�_ �_�_�_�?�_o#o5o GoYoko}o�o�o�o�o �o�o�o1CU gy�_�����_ �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q��y� ����˟�۟��%� 7�I�[�m�������� ǯٯ����!�3�E��W�i��� �$EN�ETMODE 1�U�� W ���������»��RROR_PROG %���%�����TAB_LE  ����Q�c�uσ��SEV�_NUM ��  �������_AUTO_EN�B  ̵��ݴ_;NO�� V����}��  *���������������+����(�:���FLT9R����HIS�Ð������_ALM 1]W�� �������+;����������0�?�_����  �����²u꒰T�CP_VER �!��!��@�$EX�TLOG_REQ�v������SIZ\����STK��������TOL  ���Dz~��A= ��_BWDU�*�Z�V�ǲ?�DID� ;X�Z���<��[�STEPl�~�|����OP_DO����FACTORY�_TUNv�d��D�R_GRP 1Y��`�d 	p�.°� �*u����RHB ���2 ��� �e9 ���bt �o��������J5nYA�!~}@��@�.�u��
 J��V��ȸo���_/�(/(B��  F!A�  @w�33R"�33-/@UUTn*@P  �/ȷ>u.�>*���<��ǆ-E�� F@ �"�5W�%�-J���NJk�I'P�KHu��IP��sF!���-?��  ?�/9�<�9�89�6C'6<,�5���-�V�v�7޷�t���� ��������FEAT?URE Z�V��ƱHan�dlingToo�l �5��En�glish Di�ctionary��74D St�0a�rd�6�5Anal?og I/O�7�7�gle Shif�t Outo So�ftware U�pdate%Ima�tic Back�up�9SAground Edit�0~�7Camera�0�F�?CnrRnd�ImXC�Lommo�n calib �UI�C�FnqA�@M�onitor�Kt�r�0Reliab<@�8DHCP�IZ�ata Acqu�is�CYiagn�osOA�1[ocu�ment Vie�we�BWual �Check Sa�fety�A�6ha�nced�F�:�Us�nPFr�@�7xt.� DIO �@fi�RT�Wend�PErEr�@LQR�]�Ws�Y�r�0�P E�:FCTN Menu�P�v S8gTP In�'`facNe�5Gi�gE`nrej@p Mask Exc�P�g�WHT^`Pro�xy SvoT�fi�gh-Spe�PS�ki�D�eJP�Pmm�unicN@ons�hurE`'`_�1ab�connect �2xncr``st#ru�2z>peeQP�JQU�4KAREL Cmd. L�`�ua�husRun-;Ti�PEnvkx(`�el +R@sP@S�/W�7Licen�se�Sn\�PBoo�k(System�)�:MACROs�,�b/Offse�@�uH�P8@_�pM�R�@�BP^Mech/Stop�at.p6R"�ui�RKj�x�P�0�P@)�od@wit#ch��>�EQ.����OptmЏ>��`f�iln\=�gw�uulti-T�`tC�9PCM funHw�F�o3T�R?�f�Re�gi�pr�`I�ri�gPFV����0Num� Selb����P Adju�`���J�tatu��
�iZ��5RDM Rob�ot�0scove��1F�ea7��PFreq Anly�g'Rem`��Qn�7F�>R�Servo�P��~�8SNPX b�rvNSN^`ClifQ<ɮBLibr�3鯢�0 q�����o�ptE`ssag?��4��a -C��;��/I_m>B�MILIBk�E�?P Firm6BU��PEcAcck@sKT�PTX_C�eln����F��1�V�or�qu@imulah�A�A�u��Pa�q�U�j@�Ã&�`ev�.B�.@riP޿�USB port- �@iP�PagP��?R EVNT�ϗ�nexcept�P`��t��ſX�]VC�Ar�b�bf�V2PҦ�h$����SܠSCص�V�SGEk�a�UI~�;Web Pl!� �ާ��Խ`�TeQf�ZDT Appl��d�:�ƺ� �Gri=dV�play�R�WD4�R
�.�:n�EQ�+��r-10iA/�7L*��1Grapghic���5dv�S7DCSJ�ck�q�5�larm Cau�se/��ed�8A�scii�a��LosadnP�Upl,�2�Ol�0�AGu�6N�`���yFyc@�r��0���PV��Jo��m� c�R���c���m�./�����Q�2*u:e�RAJ��P�ٶ4eqiqnL����8NRT����9On�0e He�l�HJ�`oI�alletiz?�H������_�tr�[ROS GEth�q��T@e�װ��!�n�%�2D�tP�kg&Up9g~�(2DV-�3D Tri-jQ:EAưDef.qEBa)pdei���, �bImπF�fЎ�nsp.q=�46�4MB DRAM�Z,#FRO5/@e3ll�<�Mshf!r/"�'c%3@pLƖ,ty@s˒xG��m��.[�� ��BUp���Q�B�=mai�P�߫�]Q����@q6wl!u����^`�xR�?eL� Sup������0�P�`cr��@�R����b䚮�pr1uest�rt~QQ��ߋ�L!�4O��q$�K���l Bui7�n���APLCOO�EV�l%��CGU�OCR�G�O��DR��O
TL�S_��BU/_��K��qN_d�TA�OxVB��_�W�ܑZ���_TC�B�_�V�_�W���WF +o�V�O�W._�W�ņoTEH�o�f�O�gt&�oTEj�xVF�_w�_xVGoTwBTw~o2xVH�xVIA��vL�xVLN�yUMz �bo�f_xVN�xV!P���^xVR&xV!S��܇ʏ��W���v���VGF:�L�P2_h��h�V�h��_g�D��h�FFoh���g�RD�� TUT&��01:�L�2V�L��TBGG��v�ra�in�UI��
%HsMI���pon��m�f�"�F�>&KAREL9� ��TPj��<6 SW�IMESTڢF0O�<5�
"a�X�j��� ����ͿĿֿ���'� �0�]�T�fϓϊϜ� ����������#��,� Y�P�bߏ߆ߘ��߼� ��������(�U�L� ^����������� ����$�Q�H�Z��� ~�������������  MDV�z� �����
 I@Rv��� ���///E/</ N/{/r/�/�/�/�/�/ �/???A?8?J?w? n?�?�?�?�?�?�?O �?O=O4OFOsOjO|O �O�O�O�O�O_�O_ 9_0_B_o_f_x_�_�_ �_�_�_�_�_o5o,o >okoboto�o�o�o�o �o�o�o1(:g ^p������ � �-�$�6�c�Z�l� ��������Ə���� )� �2�_�V�h����� ��������%�� .�[�R�d��������� ������!��*�W� N�`������������ ޿���&�S�J�\� �πϒϤ϶������� ��"�O�F�X߅�|� �ߠ߲��������� �K�B�T��x��� �����������G� >�P�}�t��������� ����C:L yp������ 	 ?6Hul ~�����/� /;/2/D/q/h/z/�/ �/�/�/�/?�/
?7? .?@?m?d?v?�?�?�? �?�?�?�?O3O*O<O iO`OrO�O�O�O�O�O �O�O_/_&_8_e_\_ n_�_�_�_�_�_�_�_ �_+o"o4oaoXojo|o �o�o�o�o�o�o�o' 0]Tfx�� �����#��,� Y�P�b�t��������� ������(�U�L� ^�p����������ܟ ���$�Q�H�Z�l� ~��������د���� �M�D�V�h����  H55�2}���21��R7�8��50��J61�4��ATUPͶ5�45͸6��VCA�M��CRI�UI�Fͷ28	�NREv��52��R63���SCH��DOCV�]�CSU��869zͷ0ضEIOC9��4��R69��ES�ET���J7��R{68��MASK���PRXY!�7��OCO��3帨���̸m3�J6˸53���H2�LCH��OP�LG�0�MHCuR��S{�MCS��0��55ضMDS�W���OP�MP�R�M�@�0̶PCM �R0���ض�ж@�51�51<�0n�PRS��69��FRD�FREQn��MCN��93̶�SNBAE�3�SH�LB��M��M���2�̶HTC�TMI�L����TPA��T7PTX��EL�����8������J95n,�TUT�95�wUEV��UEC��wUFR�VCC���O��VIP�CS�C,�CSG8�r�IWEB�HTTf�R6C�N�CG{IG��IPGS)�RC�DG�H7u7��6ضR85�ƷR66�R7��Rn:�R530�680�I2�q�J��H�6<�E6,�RJح�0�4��6o64\�5�N�VD��R6��R8�4Tg����8�9�0\���J93�91Đ 7+���,�D0:oF�CLI����CMS�� �ST�Y��TO�q���7v�NN�ORS�ֱJ% ��j�OL(E�ND��L��Sf(F;VR��V3D���wPBV,�APL��wAPV�CCG䶷CCR|�CD��C�DL@CSBt�C�SK��CT�CT!BL9��U0,(C��y0L8C��TC �y0�'�TC(7TC��CT1E\��07TEh��0V��TFd8F,(GL8)GI�8H�8I��E@\�87�CTM,(M�8UM@8N�8PHHPL8YRd8(TSd8W�In@VGF�GP2���P2���@�H{7VP�D�HF �VPSGVPR�&VT��YP���VTB7Vs�IHb��VI aH'VK��=VGene���� �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=?�O?a?s?�?  H55hT�1�1�[U�3R78�<50ޭ9J614�9AT�U�T�4545�<6έ9VCA�D�3CR�I,KUI8T�528n-JNRE�:52JwR63�;SCH�9/DOCV�JCU�4�869�;0�:EI�O�TsE4�:R69�JESET�;KJ�7KR68�JMA{SK�9PRXYML]7�:OCO\3�<h�J)P�<3|ZJ6�<�53�JH�\LCH^\ZOPLG�;0�Z�MHCR]ZSkMkCS�<0,[55�:�MDSW}k�[OP��[MPR�Z�@�\0n�:PCMLJR0�k�)P�:)`�[51K5u1|0JPRS[�69|ZFRD<JFwREQ�:MCN�:{93�:SNBA}K^�[SHLB�zM�{t�@ll2�:HTC�:�TMIL�<�JTP�A�JTPTX�EL�z)`�K8�;�0�JwJ95\JTUT�[�95|ZUEVZU�EC\ZUFR<JV�CC��O<jVIP�,�CSC\�CSGtlJ�@I�9WEB�:7HTT�:R6{L���CG{�IG[�IP�GS��RC,�DG��[H77�<6�:R�85�JR66JRu7[R|R53{K68|2�Z�@Jml*,|6|6\JR�\	Pj|4L�6�64���5�kNVDZR6+kR84<���IP,��8��90���KJ9&�\91��̫7[KIP�\JD0�F��CL9I�lKCMS�J9�n�:STY,�TO�:��@�K7�LNN|ZO�RS<jJ��MZZ|O]LK�END�:L��S��FVR�JV3�D,�KKPBV\�A�PL�JAPV�ZC�CG�:CCRjC�D�CDL̚CS�B�JCSK�jCTK�CTB��\���\��C�z���CL�TC�LJ�l�TC��TC�ZCTE�J��|�T�E�J��<�TF��FJ\�G��G��l�Hl��I�z)�l�k�CTM�\�M\�M��Nl�P�,�P��R��;�TSr��W��̚VGF��P2��P2�z ��VPDFLJV�P;�VPR��VT��;� �JVTB��V�KIH�VِM�<��VK,�V{�Gene�8�83EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{?��7�0STD~�4LANG�4 �9�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� ��2�D�V�RBT�6OPTNm�������� Ǐُ����!�3�E� W�i�{�������ß�5DPN�4����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}�x�ߡ߳�ted �4 �8��������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������@��ǯٯ�������*�<�N�`�r���9�9���$FEAT�_ADD ?	��������  	��ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu�����DEMO Z��?   ���} ��'��0�]�T�f� �������������� #��,�Y�P�b����� ������������ (�U�L�^��������� ���ܯ���$�Q� H�Z���~�������� ؿ��� �M�D�V� ��zόϦϰ������� �
��I�@�R��v� �ߢ߬��������� �E�<�N�{�r��� �����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo~o �o�o�o�o�o�o�o! *WN`z�� �������&� S�J�\�v��������� �ڏ���"�O�F� X�r�|�������ߟ֟ ����K�B�T�n� x�������ۯү�� ��G�>�P�j�t��� ����׿ο���� C�:�L�f�pϝϔϦ� ������	� ��?�6� H�b�lߙߐߢ����� ������;�2�D�^� h����������� ��
�7�.�@�Z�d��� �������������� 3*<V`��� �����/& 8R\����� ����+/"/4/N/ X/�/|/�/�/�/�/�/ �/�/'??0?J?T?�? x?�?�?�?�?�?�?�? #OO,OFOPO}OtO�O �O�O�O�O�O�O__ (_B_L_y_p_�_�_�_ �_�_�_�_oo$o>o Houolo~o�o�o�o�o �o�o :Dq hz������ �
��6�@�m�d�v� ������ُЏ��� �2�<�i�`�r����� ��՟̟ޟ���.� 8�e�\�n�������ѯ ȯگ����*�4�a� X�j�������ͿĿֿ ����&�0�]�T�f� �ϊϜ����������� �"�,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/
??A? 8?J?w?n?�?�?�?�? �?�?�?OO=O4OFO sOjO|O�O�O�O�O�O �O__9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿����&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t����������   ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�����y  �x�q��� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p��P����q�p�x ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p���������������$F�EAT_DEMO�IN  ��� �����IND�EX���I�LECOMP �[���B���8 SETU�P2 \B~L�  N w�5_AP2BCK� 1]B	  #�)����%����E �	���5 �Y�f��B ��x/�1/C/� g/��/�/,/�/P/�/ t/�/?�/??�/c?u? ?�?(?�?�?^?�?�? O)O�?MO�?qO O~O �O6O�OZO�O_�O%_ �OI_[_�O__�_�_ D_�_h_�_�_
o3o�_ Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0����ׯQ	� P� 2>� *.VRޯ(���*+�Q���W�{��e��PC������OFR6:��ؾg�����T   �2�����\� ��d�*.F��ϕ�	ó����qo�ߓ�STM� 9���ư%�d��ψ���HU߻�Jש�f�x���GIF�A�L��-����ߑ��JPG ����Lձ�n�����#JS�H�����6����%
JavaS�criptt���C�Se���Kֹ�v� %�Cascadi�ng Style Sheets���j�
ARGNAMOE.DT'��OЁ\;��[�k|(>k DISP*rU�Oп��� �
�TPEINS.X3ML/�:\C�cCustom Toolbar���	PASSWOR�D���FRS:�\�� %Pa�ssword Config/c�Q/ �J/�/���/:/�/�/ p/?�/)?;?�/_?�/ �??$?�?H?�?l?�? O�?7O�?[OmO�?�O  O�O�OVO�OzO_�O �OE_�Oi_�Ob_�_._ �_R_�_�_�_o�_Ao So�_woo�o*o<o�o `o�o�o�o+�oO�o s��8��n ��'���]���� �z���F�ۏj���� ��5�ďY�k������ ��B�T��x����� C�ҟg�������,��� P���������?�ί �u����(���Ͽ^� 󿂿�)ϸ�M�ܿq� ��ϧ�6���Z�l�� ��%ߴ��[����� �ߵ�D���h����� 3���W����ߍ��� @����v����/�A� ��e������*���N� ��r�����=��6 s�&��\� �'�K�o� �4�X��� #/�G/Y/�}//�/ �/B/�/f/�/�/�/1? �/U?�/N?�??�?>? �?�?t?	O�?-O?O�?�cO�?�OO(O�O�F��$FILE_DG�BCK 1]����@��� < �)
S�UMMARY.DyG�OsLMD:�O�;_@Diag� Summary�<_IJ
CONSLOG1__&Q_�_NQ�Console� log�_HK	T�PACCN�_o%�o?oJUTP A�ccountin��_IJFR6:I�PKDMP.ZI	PsowH
�o�oKU[`�Exceptio�n�oyk'PMEMCHECK5o�_*_K��QMemory� DataL�F�1l�)6qRIP�E�_$6�Zs%��q Packe�t L�_�DL�$y�	r�qSTAT����S� %~�rStatusT��	FTP���:����Vw�Qmmen�t TBD؏� �>I)ETHERNE���
q�[��NQEthern��p�Pfigura��oODDCSVRAF̏��ďݟd���� verify �all��{D�.���DIFF՟��͟xb��s��diffd���
q��CHG01 Y�@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ��VTRNDIAG.LS�̿޿s�^q=3� Ope���q� SQnostic�EWl�)VD;EV7�DATt�Q�xc�u�g�Vis��?Device�Ϫ�IMG7ºo����y�z�s�Imag�n��UP��ES��~T�FRS:\��� �OQUpdates List ��IJg�FLEXEVENQ�X�j߃�f��F� UIF E�v���B,�s��)
PSRBWLOD.CM��sL�������PPS_RO�BOWEL��GL�o�GRAPHIC�S4Dy�b�t���%4D Gra�phics Fi�leu��AOɿ��rGIG���u�
>YvGigE�ة�~�BN�? )��HADOW������\sShadow Chang���vbQRCMERR�n�\s�� CFG Er�ror�tail�� MA��C?MSGLIB� �"^o� ���T�)�ZD�����/XwZD�6 ad�HPNOTI���
/�/Zu�Notific8��H/��AGUO�/ yO?�O'?P?OOt?? �?�?9?�?]?�?O�? (O�?LO^O�?�OO�O 5O�O�OkO _�O$_6_ �OZ_�O~_�__�_C_ �_�_y_o�_2o�_?o ho�_�oo�o�oQo�o uo
�o@�odv �)�M��� ��<�N��r���� ��7�̏[������&� ��J�ُW������3� ȟڟi�����"�4�ß X��|������A�֯ e�����0���T�f� ���������O��s� �ϩ�>�Ϳb��o� ��'ϼ�K����ρ�� ��:�L���p��ϔߦ� 5���Y���}���$�� H���l�~���1��� ��g���� �2���V� ��z�	�����?���c� ��
��.��Rd�� ���M�q �<�`��� %�I��/� 8/J/�n/��/!/�/ �/W/�/{/?"?�/F? �/j?|??�?/?�?�?��$FILE_F�RSPRT  ����0�����8MDON�LY 1]�5�0� 
 �)M�D:_VDAEX?TP.ZZZ�?�?�_OnK6%N�O Back f�ile 9O�4S�6Pe?�OOO�O�?�O __?>_�Ob_t__�_ '_�_�_]_�_�_o(o �_Lo�_po�_}o�o5o �oYo�o �o$�oH Z�o~��C� g��	�2��V�� z������?�ԏ�u��
���.�@��4VIS�BCKHA&C*�.VDA�����F�R:\Z�ION\�DATA\v�����Vision VD�B��ŏ��� '�5��Y��j���� ��B�ׯ�x����1� ��үg�������X��� P��t���Ϫ�?�ο c�u�ϙ�(Ͻ�L�^� �ς��)���M���q�  ߂ߧ�6���Z���� ��%��I�������:�LUI_CONF�IG ^�5|m��� $ h�F{�5������)�;�I���|xq�s��� ��������a���  $6��Gl~�� �K��� 2 �Vhz���G ���
//./�R/ d/v/�/�/�/C/�/�/ �/??*?�/N?`?r? �?�?�???�?�?�?O O&O�?JO\OnO�O�O )O�O�O�O�O�O_�O 4_F_X_j_|_�_%_�_ �_�_�_�_o�_0oBo Tofoxo�o!o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� �����ʏ܏��� $�6�H�Z�l������ ��Ɵ؟ꟁ�� �2� D�V�h���������¯ ԯ�}�
��.�@�R� d�����������п� y���*�<�N�`��� �ϖϨϺ�����u�� �&�8�J���[߀ߒ� �߶���_������"� 4�F���j�|���� ��[�������0�B� ��f�x���������W� ����,>��b t����O���(:�  �xFS�$FL�UI_DATA �_������uRESULT 2`��� �T��/wizard�/guided/�steps/Expertb��/ /+/=/O/a/s/�/�/��*�Conti�nue with{ G�ance�/ �/�/??(?:?L?^?�p?�?�?�? T-�U��90 �`� �?���9��ps�?0OBOTOfOxO �O�O�O�O�O�O�O�  �_/_A_S_e_w_�_ �_�_�_�_�_�_n�?��?�?�<Frip �Oo�o�o�o�o�o �o�o!3E_i {������� ��/�A�S�o$on��HoAO�TimeUS/DST[� �����+�=�O�a��s������'Enabl�/˟ݟ��� %�7�I�[�m������T�?{�ݯ����Æ24Ώ3�E�W�i� {�������ÿտ翦� ���/�A�S�e�wω� �ϭϿ������ϴ�Ư�د� G��Region�χߙ߽߫� ��������)�;�+�America sou�������������)�;��?�y��#߅�G�Y��ditorL������� #5GYk}��+� Touch P�anel �� (�recommen�)���*�<N`r��U���e�w��������accesd�./@/R/d/ v/�/�/�/�/�/�/Q|�Connect� to Network�/(?:?L?^? p?�?�?�?�?�?�?�?
Y���������!/��Introducts߆O�O�O �O�O�O�O__(_:_ U^_p_�_�_�_�_�_��_�_ oo$o6oHo e�Oeo?O�X_�o �o�o�o'9K ]o��R_��� ���#�5�G�Y�k��}�����h`�ooj }oߏ�o��*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ쯫� ��Ϗ1��X�j�|��� ����Ŀֿ����� 0��A�f�xϊϜϮ� ����������,�>� ��_�!���E��߼��� ������(�:�L�^� p���߸�������  ��$�6�H�Z�l�~� ��O߱�s�������  2DVhz�� ������
. @Rdv���� ����/��'/��� `/r/�/�/�/�/�/�/ �/??&?8?�\?n? �?�?�?�?�?�?�?�? O"O4O�UO/yO�O O?�O�O�O�O�O__ 0_B_T_f_x_�_I?�_ �_�_�_�_oo,o>o Poboto�oEO�OiO�o �o�O(:L^ p�������_  ��$�6�H�Z�l�~� ������Ə؏�o�o�o �/��oV�h�z����� ��ԟ���
��.� �R�d�v��������� Я�����*���� ����C�����̿޿ ���&�8�J�\�n� ��?��϶��������� �"�4�F�X�j�|ߎ� M�_�q��ߕ����� 0�B�T�f�x���� ���������,�>� P�b�t����������� ���߱���%��L^ p�������  $��5Zl~ �������/  /2/��S/w/9�/ �/�/�/�/�/
??.? @?R?d?v?�?�/�?�? �?�?�?OO*O<ONO `OrO�OC/�Og/�O�/ �O__&_8_J_\_n_ �_�_�_�_�_�_�?�_ o"o4oFoXojo|o�o �o�o�o�o�O�o�O �O�oTfx��� ������,��_ P�b�t���������Ώ �����(��oI� m��C�����ʟܟ�  ��$�6�H�Z�l�~� =�����Ưد����  �2�D�V�h�z�9��� ]���ѿ����
��.� @�R�d�vψϚϬϾ� �Ϗ�����*�<�N� `�r߄ߖߨߺ��ߋ� տ����#��J�\�n� ������������� �"���F�X�j�|��� ������������ ������u7�� ����,> Pbt3����� ��//(/:/L/^/ p/�/ASe�/��/  ??$?6?H?Z?l?~? �?�?�?�?��?�?O  O2ODOVOhOzO�O�O �O�O�O�/�/�/_�/ @_R_d_v_�_�_�_�_ �_�_�_oo�?)oNo `oro�o�o�o�o�o�o �o&�OG	_k -_������� �"�4�F�X�j�|�� ����ď֏����� 0�B�T�f�x�7��[ �������,�>� P�b�t���������ί �����(�:�L�^� p���������ʿ��� ���џӿH�Z�l�~� �Ϣϴ����������  �߯D�V�h�zߌߞ� ����������
��ۿ =���a�s�7ߚ��� ��������*�<�N� `�r�1ߖ��������� ��&8J\n -�w�Q������ "4FXj|� �������// 0/B/T/f/x/�/�/�/ �/���/?�>? P?b?t?�?�?�?�?�? �?�?OO�:OLO^O pO�O�O�O�O�O�O�O  __�/�/�/?i_+? �_�_�_�_�_�_�_o  o2oDoVoho'O�o�o �o�o�o�o�o
. @Rdv5_G_Y_� }_����*�<�N� `�r���������yoޏ ����&�8�J�\�n� ��������ȟ��� ��4�F�X�j�|��� ����į֯����ˏ �B�T�f�x������� ��ҿ�����ٟ;� ��_�!��ϘϪϼ��� ������(�:�L�^� p߁ϔߦ߸�������  ��$�6�H�Z�l�+� ��Oϱ�s��������  �2�D�V�h�z����� ����������
. @Rdv���� }�������<N `r������ �//��8/J/\/n/ �/�/�/�/�/�/�/�/ ?�1?�U?g?+/�? �?�?�?�?�?�?OO 0OBOTOfO%/�O�O�O �O�O�O�O__,_>_ P_b_!?k?E?�_�_{? �_�_oo(o:oLo^o po�o�o�o�owO�o�o  $6HZl~ ���s_�_�_�� �_2�D�V�h�z����� ��ԏ���
��o.� @�R�d�v��������� П�������� ]����������̯ޯ ���&�8�J�\�� ��������ȿڿ��� �"�4�F�X�j�)�;� M���q��������� 0�B�T�f�xߊߜ߮� m���������,�>� P�b�t�����{� �ϟ����(�:�L�^� p���������������  ��6HZl~ ������� ��/��S�z�� �����
//./ @/R/d/u�/�/�/�/ �/�/�/??*?<?N? `?�?C�?g�?�? �?OO&O8OJO\OnO �O�O�O�Ou/�O�O�O _"_4_F_X_j_|_�_ �_�_q?�_�?�_�?�_ 0oBoTofoxo�o�o�o �o�o�o�o�O,> Pbt����� ����_%��_I�[� ��������ʏ܏�  ��$�6�H�Z�~� ������Ɵ؟����  �2�D�V��_�9��� ��o�ԯ���
��.� @�R�d�v�������k� п�����*�<�N� `�rτϖϨ�g����� ������&�8�J�\�n� �ߒߤ߶��������� ��"�4�F�X�j�|�� �������������� ����Q��x������� ��������,> P�t����� ��(:L^ �/�A��e����  //$/6/H/Z/l/~/ �/�/a�/�/�/�/?  ?2?D?V?h?z?�?�? �?o���?�O.O @OROdOvO�O�O�O�O �O�O�O�/_*_<_N_ `_r_�_�_�_�_�_�_ �_o�?#o�?Go	Ono �o�o�o�o�o�o�o�o "4FXio|� �������� 0�B�T�ou�7o��[o ��ҏ�����,�>� P�b�t�������iΟ �����(�:�L�^� p�������e�ǯ��� ����$�6�H�Z�l�~� ������ƿؿ�����  �2�D�V�h�zόϞ� ���������Ϸ��ۯ =�O��v߈ߚ߬߾� ��������*�<�N� �r��������� ����&�8�J�	�S� -�w���c��������� "4FXj|� �_����� 0BTfx��[� �������/,/>/ P/b/t/�/�/�/�/�/ �/�/�?(?:?L?^? p?�?�?�?�?�?�?�? ����EO/lO~O �O�O�O�O�O�O�O_  _2_D_?h_z_�_�_ �_�_�_�_�_
oo.o @oRoO#O5O�oYO�o �o�o�o*<N `r��U_��� ���&�8�J�\�n� ������couo�o鏫o �"�4�F�X�j�|��� ����ğ֟蟧��� 0�B�T�f�x������� ��ү������ُ;� ��b�t���������ο ����(�:�L�]� pςϔϦϸ�������  ��$�6�H��i�+� ��O������������  �2�D�V�h�z��� ]���������
��.� @�R�d�v�����Y߻� }����ߣ�*<N `r������ ���&8J\n ��������� /��1/C/j/|/�/ �/�/�/�/�/�/?? 0?B?f?x?�?�?�? �?�?�?�?OO,O>O �G/!/kO�OW/�O�O �O�O__(_:_L_^_ p_�_�_S?�_�_�_�_  oo$o6oHoZolo~o �oOO�OsO�o�o�O  2DVhz�� �����_
��.� @�R�d�v��������� Џ⏡o�o�o�o9��o `�r���������̟ޟ ���&�8��\�n� ��������ȯگ��� �"�4�F���)��� M���Ŀֿ����� 0�B�T�f�xϊ�I��� ����������,�>� P�b�t߆ߘ�W�i�{� �ߟ���(�:�L�^� p���������� ���$�6�H�Z�l�~� �������������� ��/��Vhz�� �����
. @Qdv���� ���//*/</�� ]/�/C�/�/�/�/ �/??&?8?J?\?n? �?�?Q�?�?�?�?�? O"O4OFOXOjO|O�O M/�Oq/�O�/�O__ 0_B_T_f_x_�_�_�_ �_�_�_�?oo,o>o Poboto�o�o�o�o�o �o�O�O%7�_^ p�������  ��$�6��_Z�l�~� ������Ə؏����  �2��o;_���K ��ԟ���
��.� @�R�d�v���G����� Я�����*�<�N� `�r���C���g���ۿ ����&�8�J�\�n� �ϒϤ϶����ϙ��� �"�4�F�X�j�|ߎ� �߲����ߕ�����˿ -��T�f�x���� ����������,��� P�b�t����������� ����(:��� �A�����  $6HZl~ =�������/  /2/D/V/h/z/�/K ]o�/��/
??.? @?R?d?v?�?�?�?�? �?��?OO*O<ONO `OrO�O�O�O�O�O�O �/�O�/#_�/J_\_n_ �_�_�_�_�_�_�_�_ o"o4oE_Xojo|o�o �o�o�o�o�o�o 0�OQ_u7_�� ������,�>� P�b�t���Eo����Ώ �����(�:�L�^� p���A��eǟ���  ��$�6�H�Z�l�~� ������Ưد�����  �2�D�V�h�z����� ��¿Կ�������+� �R�d�vψϚϬϾ� ��������*��N� `�r߄ߖߨߺ����� ����&��/�	�S� }�?Ϥ���������� �"�4�F�X�j�|�;� ������������ 0BTfx7��[� �����,> Pbt����� ���//(/:/L/^/ p/�/�/�/�/�/�� ��!?�H?Z?l?~? �?�?�?�?�?�?�?O  O�DOVOhOzO�O�O �O�O�O�O�O
__._ �/�/?s_5?�_�_�_ �_�_�_oo*o<oNo `oro1O�o�o�o�o�o �o&8J\n �?_Q_c_��_�� �"�4�F�X�j�|��� ����ď�oՏ���� 0�B�T�f�x������� ��ҟ����>� P�b�t���������ί ����(�9�L�^� p���������ʿܿ�  ��$��E��i�+� �Ϣϴ����������  �2�D�V�h�z�9��� ����������
��.� @�R�d�v�5ϗ�Yϻ� }������*�<�N� `�r������������� ��&8J\n ���������� ��FXj|� ������// ��B/T/f/x/�/�/�/ �/�/�/�/??�# �G?q?3�?�?�?�? �?�?OO(O:OLO^O pO//�O�O�O�O�O�O  __$_6_H_Z_l_+? u?O?�_�_�?�_�_o  o2oDoVohozo�o�o �o�o�O�o�o
. @Rdv���� }_�_�_�_��_<�N� `�r���������̏ޏ �����o8�J�\�n� ��������ȟڟ��� �"����g�)��� ����į֯����� 0�B�T�f�%������� ��ҿ�����,�>� P�b�t�3�E�W���{� ������(�:�L�^� p߂ߔߦ߸�w�����  ��$�6�H�Z�l�~� ����������� ��2�D�V�h�z����� ����������
-� @Rdv���� �����9�� ]������� �//&/8/J/\/n/ -�/�/�/�/�/�/�/ ?"?4?F?X?j?)�? M�?qs?�?�?OO 0OBOTOfOxO�O�O�O �O/�O�O__,_>_ P_b_t_�_�_�_�_{? �_�?oo�O:oLo^o po�o�o�o�o�o�o�o  �O6HZl~ �������� �_o�_;�e�'o���� ��ԏ���
��.� @�R�d�#�������� П�����*�<�N� `��i�C�����y�ޯ ���&�8�J�\�n� ��������u�ڿ��� �"�4�F�X�j�|ώ� �ϲ�q�������	�˯ 0�B�T�f�xߊߜ߮� ���������ǿ,�>� P�b�t������� ������������[� ߂�������������  $6HZ�~ �������  2DVh'�9�K� �o����
//./ @/R/d/v/�/�/�/k �/�/�/??*?<?N? `?r?�?�?�?�?y�? ��?�&O8OJO\OnO �O�O�O�O�O�O�O�O _!O4_F_X_j_|_�_ �_�_�_�_�_�_o�? -o�?QoOxo�o�o�o �o�o�o�o,> Pb!_����� ����(�:�L�^� o�Ao��eog�܏�  ��$�6�H�Z�l�~� ������s؟����  �2�D�V�h�z����� ��o�ѯ�����˟.� @�R�d�v��������� п����ş*�<�N� `�rτϖϨϺ����� �������/�Y�� �ߒߤ߶��������� �"�4�F�X��|�� ������������� 0�B�T��]�7߁��� m�������,> Pbt���i�� ��(:L^ p���e�w����� ���$/6/H/Z/l/~/ �/�/�/�/�/�/�/�  ?2?D?V?h?z?�?�? �?�?�?�?�?
O�� �OO/vO�O�O�O�O �O�O�O__*_<_N_ ?r_�_�_�_�_�_�_ �_oo&o8oJo\oO -O?O�ocO�o�o�o�o "4FXj|� �__������ 0�B�T�f�x������� moϏ�o�o�,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ���!��E��l�~� ������ƿؿ����  �2�D�V��zόϞ� ����������
��.� @�R��s�5���Y�[� ��������*�<�N� `�r����g����� ����&�8�J�\�n� ������c��������� ��"4FXj|� �������� 0BTfx��� ����������#/ M/t/�/�/�/�/�/ �/�/??(?:?L? p?�?�?�?�?�?�?�?  OO$O6OHO/Q/+/ uO�Oa/�O�O�O�O_  _2_D_V_h_z_�_�_ ]?�_�_�_�_
oo.o @oRodovo�o�oYOkO }O�O�o�O*<N `r������ ��_�&�8�J�\�n� ��������ȏڏ��� �o�o�oC�j�|��� ����ğ֟����� 0�B��f�x������� ��ү�����,�>��P��!�3������$�FMR2_GRP� 1a���� �C4 w B�[�	 [��߿�ܰE�� �F@ 5W��S�ܰJ��NJ�k�I'PKH�u��IP�sF�!���?�  �W�S�ܰ9�<9��896�C'6<,5����A�  l�Ϲ�BHٳB�հ�����@�33�33S�۴��ܰ/@UUT'�@��8���W�>u.�>*���<����=�[�B=���=�|	<�K�<�q�=�mo����8�x	7�H<8�^6�Hc7��x?� ���������"��F��X���_CFG =b»T Q������X�NO ^º
F0�� ���W�RM_CHKTYP  ��[�ʰ�̰����ROM�_�MIN�[����9����X��SSB�h�c�� ݶf�[�]�����^�TP_DEF_�O�[�ʳ��I�RCOM���$�GENOVRD_�DO.�d���TH�R.� dd��_�ENB�� ��RWAVC��dO�Z�� ���Fs  �G!� GɃ��I�C�I(i J���+���%�q���� �Q�OU��j¼��8����<6�i��C�;]�[�C�  D�+��3@���B���p�.��R SMT���k_	ΰ\��$HoOSTCh�1l¹�[��d�۰ M5C[���/Z�  27.0� =1�/  e�/? ?'?9?G:�/j?|?�?�?�,Z?T3	anonymouy �?�?�	OO-O?N�/ڰRH RK�/�?�O�/�O�O�O �O_V?3_E_W_i_�O &_�?�_�_�_�_�_@O �_dOvOSo�_�Ojo�o �o�o�o_�o+ =`o�_�_���� �o&o8oJoL9��o ]�o��������oɏۏ ����4�j+�Y�k� }��������� � �T�1�C�U�g����� ������ӯ��x�>�� -�?�Q�c�����Ο�� �Ͽ����)�;� ��_�qσϕϧ�ʿ � �����%�7�~��� ��߶ϣ�������� ���Ϻ�3�E�W�i�� ���ϱ���������@� R�d�v�x�J��߉��� ���������+ =`���������:$h!ENT 1=m P!V  7 ?. c&�J�n�� �/�)/�M//q/ 4/�/X/j/�/�/�/�/ ?�/7?�/?m?0?�? T?�?x?�?�?�?O�? 3O�?WOO{O>O�ObO �O�O�O�O�O_�OA_ _e_(_:_�_^_�_�_��_�ZQUICCA0�_�_�_?od1@oo.o�od2�olo~o��o!ROUTE�R�o�o�o/!P�CJOG0!�192.168�.0.10	o�SC�AMPRT�\!�pu1yp��vRT��o��� !S�oftware �Operator? Panel�m�n��NAME �!�
!ROBO��v�S_CFG �1l�	 ��Auto-s�tarted'�FTP2��I�K 2��V�h�z������� ԟ����	���@� R�d�v���	����� ��:���)�;�M�_� &���������˿�p� ��%�7�I�[��"� 4�F�ڿ�������� !�3���W�i�{ߍߟ� ��D���������/� vψϚ�w�ߛ��Ͽ� ��������+�=�O� a�������������� ��8�J�\�n�p�]�� ��������� #5X�k}� ���0/D 1/xU/g/y/�/RH/ �/�/�/�//?�/?? Q?c?u?�?���/ ?�?:/O)O;OMO_O &?�O�O�O�O�O�?pO __%_7_I_[_�?�? �?t_�O�_O�_�_o !o3o�OWoio{o�o�_ �oDo�o�o�o�����_ERR n���-=vPDUSI�Z  �`^�P��Tt>muWRD �?΅�Q�  �guest �f������~��SCDMNGRPw 2o΅Wp���Q�`���fK�L� 	P01.�05 8�Q  � �|��  �;|��  ~z[ ���w����*���Ť�x����[ݏȏ���בPԠ�������)����D�r���؊p"*�Pl�P���Dx���dx�*�����%�_GWROU7�pLyN���	/�o���QU%P��UTu� ��TYàL}?pT�TP_AUTH �1qL{ <!iPendan���o֢!KAREL:*�������KC��ɯۯ���VISION SET�9����P�>� h��f�����������ҿ����X�CTRL rL}O�u���a
��pFF�F9E3-ϝTF�RS:DEFAU�LT��FAN�UC Web Server�ʅ�t� X���t@���1�C��U�g�;tWR_CONFIG s;�� ��=qIDL_CPU_PC����aBȠP�� BH��MIN�܅q��?GNR_IOFq{r��`Rx��NPT_S_IM_DO���STAL_SCR�N� �.�INT�PMODNTOL8Q����RTY0���8�-�\�ENBQ�-����OLNK 1tL{�p�������)�;�M���MAST�E�%���SLAV�E uL|�RA?MCACHEk�c�}O^�O_CFG�������UOC�����CMT_OP���Pz�YCL������_?ASG 1v;��q
 O�r��� ����&8pJ\W�ENUMzs5Py
��IP����RTRY_CN���M�=�zs���Tu ������w���p/��p��P_MEMB?ERS 2x;�l�k $��X"��?��Q'W/i)��RCA_�ACC 2y��  Y�h k�%�� 6��" � !pQ�`�&4�@�p@�/�&s��$�(��$BUF001 �2z�= �Z�u0  u0�k�:4z:4�:4�:4��:4�:4�:4�:4�Z:4�:3��4 �4U/�4A�4P�4a�4Uq�4��4��4��4U��4Ċ4Ԋ4�4��:3�DD'�D6DGDWDh�DrJ�  JЭ�Y4��JD�JD�jJD�JD�:3�rDUrD"rD1rDCrDURrDdrDtrD�rDU�rD�rD�rD�rDU�rD�rD�:4	:4U:4*:49:4J:392$?63:1@1ERI0 ERQ0ERY0ERa0ERi0 ERq0ERy0ER�0ER�0 :1�1�R�0�R�0�R�0 �R�0�R�0�R�0�R�0 �R�0�R�0�R�0�R�0 �R�0�R�0�R@:1A b@b@b!@b)@ b1@b9@bA@BAHO?u0`�@`A:1 hAmbq@:1xA}b�@}b �@}b�@}b�@}b�@}b �@}b�@}b�@}b�@}b �@}b�@}b�@}b�@}b �@}b�@ER�@ERPER�	PERPERP:193 -_65GSNrI2WSVrY2 gSVri2wSVry2�SVr �2�S�r�2�S�r�2�S �r�2�S�r�2�S�r�2 �S�r�2�S�r�2c�� Cc�B'c�)B7c �9BGc��QcO`QBO` YBO`aBocV�qBc�� �B�c���B�c���B�c ���B�c���B�c���B �c���B�c���B�cVr RsVrRs�Ԝ!��2{�4r�}ŋ���<����o�o��2��HIS!2}� �ܷ! 2024O-08-"0����П�����'��  3 ���o�� �m�Q�c���X�RX��7-25�������Ư���� 7 ;RXj�4 ӯ�p�*�<�s��cȅ��O���������ܩ  �;�´`t�" *c� N���������t��bꅨ2 m�Z�l�~ϐϻ�Ѱm�b�K���������}���fn��6-27�I�6�H�Zߵ�ǺĲf�n�Ϥ߶�����}��g�6%��$�6�`m�o�ɲo���g��������}��j�@ؐ������ح�1��J�űj�óX� j�|���q��,P���� ������#5G5��� +A�o�d� : M ��y�y��������1�9� _�8 �+=OaO�a������ߦ,r�JDɰV�cѰ�ٰ:j �/)/;/)�;ϖ�/P�/�/�/��;L�b�� i�/�/??��r/@_?q?�?ݨ��d�d���/�?�?�? O��  �6OHOZOحiɰi �5m�?�O�O�O�O��@�_$_6_�?�3:�! �5J��2Q�2D_�_�_ �_��3r����_o$o 6oHoZolo5�" aA� �bn �b�o�o��o�o�!�a�o K]o����o����ګ�b�Ѱ �qٰ�*�<�N�`�N/�`/�����̏ޏ�� ��������*�<�*? <?��������ݨ��ɰ ����������%� O%O[�m����ȟl� ޟ˯ݯ���O�o7�I�[�H��~�Ѱ~� I���Q𺯯���ӿ�_�A_I_CFG �2~�[ H
�Cycle Ti�me(�Bus}y�Idl�N-�mi���S��Up� �R�ead(�Do�wG�C�r X��C�ount �	Num �.�����(�y����PROG����U�P�)�/softpar�t/genlin�k?curren�t=menupa�ge,1133,��W:�L�^�p�K̤�S�DT_ISOLCw  �Y� ����J23_DSP_ENB  ���T���INC ����(���A   ?�^ =���<#��
���:�o ��2�D�(�/�l���OB��C��O��ֆ��G_GROUP �1���i< �������t�E?����(�Q'� L�^�p�/�����������\�~�G_IN�_AUTO����P�OSRE���KA�NJI_MASK�0��DRELMO�N ��[��(�y ��������fJ�Ã����(�|-��KCL_L �NUM��G$KE�YLOGGING�D�P�zQ����LA�NGUAGE ��U��DEFAULT �6�QLG�����S���(�x�  {8T�H  �(�K'0縤(�qQ�ލ�;��
*!(�UT1:\ J/ L/Y/k/}/�/�/�/ �/�/�/�/$>(�H?��VLN_DISP ���P�&�$�^4�OCTOL|�Dz�����
�1GBOOK ��}Q1V�11}P�@*O!O 3OEOWOiKyM�TËIgF	�5)����O�}���2_BUFF� 2��� �O��_|R��6_M� R_d_�_�_�_�_�_�_ �_�_o3o*o<oNo`o��o�o�o�o���ADCS ������L �O��+=Oa�d�IO 2��k !������� ������*�:� L�^�r���������ʏ ܏���$�6�J�uu�ER_ITM��d ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����7x��SEVD��t�TYP����s�������)RSTe�eS�CRN_FL 2��}������/�A�S�e�wϨ�TP�{��b��=NGN�AM��E��dUPMSf0GI��2��}��_LOAD���G %��%D�ROP_�EIT�O_3�ϑ�MAXUALRMb2�@����
K���_P�R��2  �3�AK�Ci0��qO=_'X��ެ�P 2��; ��*V	����
*����4��*��'� `�	xN��z���� �������1�C�&�g� R���n����������� 	��?*cFX ������� ;0q\�� �����/�/ I/4/m/X/�/�/�/�/ �/�/�/�/!??E?0? i?{?^?�?�?�?�?�? �?�?OOAOSO6OwO�bO�OD�DBG*� ���գѢѤO�@_LDXDISA�����ssMEMO_A�P��E ?��
 �Ax$_6_H_�Z_l_~_�_�_K�FR�Q_CFG �ږ��CA w@�4�S�@<��d%�\o�_�P�Ґ��^��*Z`/\b **:eb�DXojh o�F�o�o�o�o�o �o;�O��dZ�U0�y|��z,(9� Mt���1��B�g� N���r��������̏�	���?�A�ISCg 1���K` ��O �����O���O֟�����K�]�_MSTR ��3��SCD 1�]��l�� {�����دïկ��� 2��V�A�z�e����� ��Կ�������@� +�=�v�aϚυϾϩ� ��������<�'�`� K߄�oߨߓߥ����� ���&��J�5�Z�� k����������� ���F�1�j�U���y� ������������0`T?x�MK�Q��,��Q�$MLoTARM�R�?g� ~s�@�|��@METPU�@�l��4�NDSP_ADCOL<�@!CMNT7(�FNSWiSTL�Ix *%� �,����Q��*_POSCF���PRPMV�STv51�,� 4�R#�
g!|qg%w/�' c/�/�/�/�/�/�/? �/?G?)?;?}?_?q?��?�?�?�?�1*SI�NG_CHK  }{$MODA�S��e���#EDE�V 	�J	M�C:WLHSIZE��Ml �#ETASK� %�J%$12�3456789 ��O�E!GTRIG ;1�,� l�Eo�#_�y_S_�}�FYP�A�u9D"CEM_�INF 1�?k�`)AT&F�V0E0X_�])��QE0V1&A3�&B1&D2&S0&C1S0=�])ATZ�_#o
d�H'oOo�QC_wohA�o�obo�o�o�o  �_&�_�_�_o�3o ��o���o��"� 4��X���AS e֏���C�0�� �f�!���q�����s� 䟗�����͏>��b� ��s���K���w��� ٯ�ɟ۟L����#� ����Y�ʿ���� $�߿H�/�l�~�1��� U�g�y����ϯ� �2� i�V�	�z�5ߋ߰ߗ�|��PONITOR��G ?kK   	EXEC1o��2�3�4�5���@�7�8�9o����(� ��4��@��L��X �d��p��|��2���2��2��2��2���2��2��2��2���2��3��3��3�(�#AR_GRP_�SV 1��[ �(�1?Ý����{b?7N���b��=.3IRM�A_DsҔN~��ION_DB-@��1Ml  ��l �FH"�+�0l �����N BL"}FI-ud1}E���)PL_N�AME !�E�� �!Defa�ult Pers�onality �(from FD�)b*RR2�� �1�L�XL��p�X  d �-?Qcu�� �����//)/ ;/M/_/q/�/�/�/f2)�/�/�/??,? >?P?b?t?f<�/�? �?�?�?�?�?
OO.O @OROdOc	�6�?�N
�O�OfP�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�_�_�O�O 2oDoVohozo�o�o�o �o�o�o�o
.@ o!ov����� ����*�<�N�`��r����� Fs�  GT�G�#Me��x �ÏՍfd�������(� 6������
 �m�~�h����� ������ ğ֟�����:���
�h]�m�f��	`��𠯲�į��:�o�Ab	����� A�  /���P� ���r�������^�˿@ݿȿ��%��R�� 1��	X ��?, � ��� ~a� @D�  t�?�z�`�?f |�f�A/��t�{	��;��	l��	 �xJ������ �� �u<�@���� ������K�K ���K=*�J����J���J9���
�ԏC߷�@�t�@{S�\҇�(Ehє��.��I���ڌ���T;f�ґ�$���3��´  ��@��>�Թ�$� � >����ӧ=Uf��x`���� �
���Ǌ���� �  {�  @T�����/  �H �l�����-�	'� �� ��I� ��  �<�+�:��È��È=��Q���0Ӂ��N �[�?�n @���f���f�k���,�<av�  '��Y����@2��@�0c@�Ш���C��}Cb C��\C�������G�@�������� )�B�b $/�!��L��Dz�o�ߓ~���0��( �� -���������!���D�  ���恀?�ff0G�*<� }�qD�1�8����>��Hbp��(�(���P���	������>�?�՚��x���W�<
�6b<߈;����<�ê<�?��<�^��I/2��A�{��fÌ¾,�?fff?_�?y&� T�@�.�"�J<?�\��"N\�5���!��(� |��/z��/j'��[0? ?T???x?c?�?�?�?`�?�?�?5��%F� �?2O�?VO�/wO�)IO��OEHG@ G@�0��G�� G} ଙO�O�O_	_B_-_\f_Q_BL��B��Aw_[_�_b��_�[�_ ��mO3o�OZo�_~o�ox�o�o���b��PV( @|po	lo- *cU�ߡA���r5eCP�Lo�}?����#���5��W�s��6�Cv�q�CH3� j�t�����q�����|^(�hA� �AL�ffA]��?��$�?��;����u�æ�)��	ff��C��#�
���g\)��"�33C�
������<��؎G�B����L�B�s?����	";��H�ۚG��!�G��WIY�E���C�+��8�I۪I�5��HgMG��3E��RC�j�=x�
�pI����G��fIV=�E<YD�C <�ݟȟ����7�"� [�F��j�������ٯ į���!��E�0�i� T�f�����ÿ���ҿ ����A�,�e�Pω� tϭϘ��ϼ������ +��O�:�s�^߃ߩ� ���߸������ �9� $�6�o�Z��~��� ���������5� �Y� D�}�h�����������@����
C.(�g���/"���<��t��q�3�8����q4�Mgu���q�V�wQ�
4p�+4�]$$dR��v���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/��/�/�/�/  %� �/�/+??O?:?s?/`�_�?�?�?�;�?��?O�? OFO4O�r LO^O�O�O�O�O�O�J  2 Fs�w�GT�V�M��uBO�|r�pp�C��S@�R_�poy_�_؝_�_o \!�WɃh_oo(o�z�?���@@�zJ�D�p�pk1�p�~
 6o�o�o �o�o�o�o);�M_q�ڊsa �����D��$�MR_CABLE� 2�� )]��T�LaMaa?�PMaLb�p�Z�ɴ&P�C�p�!O4�>�B����"��>� F�ڈ�F��"��v�_l  ��&P�v�^wdN�{0�_��V��R3���F�[�7�I�X�T��6P� C$��Č���y�2�� j&����F.S�,���| ��&Pr��C���=�����$��� Z�RK�{F�h څ��s9�"T�p�� J�D�V�h�z�ߟڟ�� ��ԟ�K�
��F�@��R�d��	j��!� ��j��������;j������@��������� �� ��`�%�j�;j*** �sOM ���y���{�  / j���%% 23456�78901ɿ۵ �ƿ���� �� AQ�� �!
�z��not sent� ���W��TESTFECS7ALG� eg�ZAQ�d��ga%�
���@���$�r�̹�������� 9UD1�:\mainte�nances.x�mS�.�@�vj��DEFAULT��\�rGRP 2���  p�R�I�%�  �%1st� mechani�cal chec�k��!���������E��Z�(��:�L�^��"��controller�����߰��D�����0 ��$�s�M��L��""8b���v��B�����������/�AC}�a�6����@dv���s�C���ge��. battery�&��E	S(:L^p�	�|�duiz�ablet  D�а���ѿ�E��/�"/4/s��gre�as��'f�r#-� |!�/�E��/�/��/�/�/s�
�oi0,�g/y/�/�/t? �?�?�?�?s��
�XֈW��1<X�AO�E
c?8OJO\OnO�OB�t��?O��'O��O_ _2_D_s�O?verhauE��L��R xXЌQ�_���O�_�_�_�_oX�$�_0oϤFi4oV� �_�o�o�o�o�oo�o @oRodo%K]o� ��o�*�� #�5�G��X�}���� �ŏ׏����\�1� C���g����������� ӟ"���F�X�-�|�Q� c�u�����蟽��� �B��)�;�M�_��� ��ү䯹��ݿ�� �%�t�IϘ����ο �ϵ�������:��^� pςϔ�i�{ߍߟ߱�  ���$�6�H�	�/�A� S�e�w��ߛ������ ������+�z�<�a� ��d������������ @�'v�K��o� ����*< `5GYk}�� ��&�//1/ C/�g/���/��/ �/�/�/	?X/-?|/�/ c?�/�?�?�?�?�?? �?B?T?f?x?MO_OqO �O�O�?�OOO,O�O _%_7_I_[_�O_�O �O�O�_�_�_�_o!o�T	 T"oOoaoso �_�o�_�k�o�o�o�o �o�o2Dz� �`r����� .�@���v�����\��n�Џ⏤����R� ��Q?�  @�a �oW�i�{���fC�����̟aX*�**  ����� � �2�D��h�z��������_�S��� ���կ7�I�[��� ��ɯ/���ǿٿ#�� �!�3�}�����{ύ� ���s�������C�U� g��S�e�w�9ߛ߭�п�	�߉e�a�$�MR_HIST �2����� 
� \jR$ 2345678901*�(2����)�9c_�� ��R��a_������� ��=�O�a��*�x��� ��r�������9 ��]o&�J�� ���#�G��k}4��d�SK�CFMAP  .��������`��ONR�EL  �����лEXCFE�NB'
��!F�NC$/$JOGO/VLIM'd�m ��KEY'p%y%_PAN(�"�"��RUN`,p%��SFSPDTY�PD(%�SIGN|/$T1MOTb/�!�_CE_G�RP 1��� �"�:`��n?�c[?�? �؆?�?~?�?�?�?!O �?EO�?:O{O2O�O�O hO�O�O�O_�O/_�O (_e__�_�_�_�_v_��_�_�_o�׻QZ_EDIT4��#�TCOM_CFG 1��'%to�o��o 
Ua_ARC�_!"��O)T_M�N_MODE6=�Lj_SPL�o2&UAP_CPL�o�3$NOCHECK� ?� � Rdv��� ������*�<��N�`��NO_WA�IT_L 7Jg50N�T]a���U	�޲�_ERR?12���ф��	��-�����R�d����`O�����| k%
aB�����o����C�������,V9<� �� ?�Uϟ�j����قPARAuMႳ��N��oR�=��o��� = e������گ� ȯ��"�4��X�j�F�<�蜿��A�ҿ�"?ODRDSP�c6�/(OFFSET_�CAR@`�o�DI�S��S_A�`A�RK7KiOPEN_FILE4�1�a�Kf�`OPTION�_IO�/�!��M_�PRG %�%c$*����h�WOT�[�E7O���8�Z��  �O�r"�÷"�	 �V�"��Z��RG�_DSBL  ���ˊ���RI_ENTTO Z�C���A �U^�`IM_D����O��V�LCT ���Gbԛa�Z=d��_PEX�`7�n*�RAT�g d/%�*��UP ���{��������|�����$PAL��������_POS_CCHU�7����2>3��L�XL�p��$�ÿU� g�y������������� ��	-?Qcu ����Y2C�� �"4FXj| ������ / /$/6/H/Z/l/~/�Y���.��/�/ςP�/??,?>?P?b? t?�?�?�?�?�?�?�? OO�/�/LO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_)O;O�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�_�<���o�m ��� ~BPw�m�m���~�jw#Ьw� �����2�T��p`��w���H��t	`��̏ޏ��:�o������ �2��pA�  I��j�`��� ������џ����@��#�)�Or�1������ 8���, ��\Ԡ�� @D��  ��?���~�?8� ���!D�������%G�  ;�	l���	 �xoJ젌������ �<� ���� ��2�H(���H3k7HS�M5G�22G�?��GN�3%�Rذ�oR�d�2�Cf��a���{�ׄ�����/��o3��¸��4���>���К�����3�A�q½{q�!�ª��ֱ� �"�(«�=�2����� ���{  @��Њ���  ���Њ�2���.�	'�� � ��I�� �  �<V�,�=�������|�ß���  �y�?�n @"��]�<߼+������-�9N�Д�  '�Ь��w�ӰC��C��\C߰��Ϲ��ߤ!��/�@�4���/�	�2�~�B��B�I�;�)�j客z+���쿱����������( �� -���#�������!��]�9��  q�?��ffaH�Z��� ��������8� ����!>�|P��}�(� ���P�������\�?W��� x� ����<
6b<߈�;܍�<�ê�<���<�^��*�gv�A)ۙ�������F�?fff?�}�?&� ��@�.���J<?�\��N\��)� ����������ޤ y�N9r]��� ����/&/�J/ 5/n/�	g/�/c(G@ G@0i�?G�� G}���/ ??<?'?`?K?�?o?WBLi�B��A�? y?�?|��?K�?ů�/ QO�/xO�?�O�O�O�O�m��b��n�t @|�O'_�OK_6_H_�_lS��A��RS�i��Cn_�_j_0O�]?Ƀ�ooAo,o¹�mWi���ToC��F�`CHQo>Jd�`�a�a@Iܚ>(�hA� �AL�ffA]��?��$�?���ź���u�æ�)��	ff��C��#�
�opg\)���33C�
������<���nG�B����L�B�s?����	0ź�H�ۚG��!�G��WIY�E���C�+��½I۪I�5��HgMG��3E��RC�j�=�~
�pI����G��fIV=�E<YD�# Zo���
��U�@� y�d���������я�� ���?�*�c�N��� r��������̟�� )��9�_�J���n��� ��˯���گ�%�� I�4�m�X���|���ǿ ���ֿ���3��W� B�Tύ�xϱϜ����� ����	�/��S�>�w� bߛ߆߿ߪ߼�����@��=�(�a�L�(qg��)����Z������a�3�8������a4�Mgu�����a�V�wQ�(�4p�+4�]B�B���p�����������UPbP���QO%x�1[FjR��������  C�� �I4mX�8`
O�������.//>/d/R/�R j/|/�/�/�/�/�/:  2 Fs�g�GT�&6�M��eBmp�R�P�aC��3@�_p?�?�?�?�?�?�=�S�OO)O�;OMO�c?���@U@�j��`�`��1�`�^
  TO�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�j�A ����D���$PARAM�_MENU ?�B�� � DEFP�ULSE{	W�AITTMOUT�kRCVo �SHELL_W�RK.$CUR_oSTYL`Dl�OPTZ1ZoPTB�ooibC?oR_DECSN`���l�o�o �o&OJ\�n������QS�SREL_ID � >�
1��uUS�E_PROG �%�Z%�@��sCC�R` �
1�SS�_H�OST !�Z!X���M�T _����x������L�_TGIMEb �h��P?GDEBUG�p�[��sGINP_FL'MSK�E�T� V��G�PGAr� 5���?��CHS�D�TY+PE�\�0�� 
�3�.�@�R�{�v��� ��ï��Я���� *�S�N�`�r������� ���޿��+�&�8πJ�s�nπϒϻ�G�W�ORD ?	�[
? 	PR2���MAI�`�SU�a��TEԀ���s	Sd�COL�h�C߸�L� C�՜~�h�d*�TR�ACECTL 1�B��Q ��� '���0�ށ�DT Q��B��М�D ȿ � �@��й��ҥ@����
�����1�@�؍@⨐��/Y ��Y��A�U	@�
@�@�@� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=?@O?a?s?�?�?�3�4� ��2�4�Y�Y� �4�4�4 ����4�(O:OLO^OpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����� ����*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟڟ���� "�4�F�P�$Or����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~�f��� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo�xo�o�o�o�o�o�a��$PGTRACE�LEN  �a � ����`��f_UP _����q'p�q p�a_CFoG �u	s�a0q�Lt�ceqx>c}  �qu4r�DEFSPD e�?|�ap��`�H_CONFIG� �us ��`�`d�t��b 	�a�qP�tcq��`ۂ�`IN7pTROL �?}_q8�u��PE�u��w��qLt�qqv�`L�ID8s�?}	v�L�LB 1��y ���B�pB4Ńqv �އ؏�	�s << �a?��'��� A�o�U�w�������۟ ��ӟ��#�	�+�Y�v�񂍯����ï
���������/�u�GRP� 1ƪ��a@�j��hs�a�A�
D�� �D@� Cŀ @�٭^�t������q�p���.� ����Ⱦ´���ʻB �)�	���?�)�c���a>��>�,᷁Ϻ��ζ� =4?9X=H�9��
� ���@�+�d�O���s���o߼�����  Dz���`
��8��� H�n�Y��}����� ��������4��X�C��|���)��
V7�.10beta1�Xv A���ι��!�����?!�G�>\=y��#��{33A!���@��͵���8wA��@�/ A�s�@Ls���� ��"4FXLs�ApLry�ā���_��@l��@W�33q�`s��k��Anff�a���ھ��)7�x�� �ar� T�n�t����	�t�KNOW_M � |uGvz�SV ��z�r�&� ���>/�/G/��a��y�MM���{� ���	^r�` (l+/�/',�$�@XLs	����@���%�"�4�.N�z�MRM��|-TU�y�c?u;e�OADBANFW�D~x�STM�1 �1�y�4Garra_B�2Sem��?~s�;Co�2��O�7��3Antena�_Full @� �VODe�qH��^OpO �O�O�O�O�O�O!_ _ _W_6_H_�_l_~_�_��b�72�<�!4�_ � �<�_�_N�3 �_�_
oo�749oKo]ooo�75�o�o�o�o��76�o�o�77 2DVh�78��X���7MA�0���swwOVLD � �{�/a�2P�ARNUM  p�;]��u�SCH*� 8�
����ω�3�UPD��[�ܵ+�>wu_CMP_r -���0�'�5C�ER�_CHKQ���`�1�"e�N�`�RS>0��?G�_MO�?_���#u_RES_G
�0��{
Ϳ@�3� d�W���{�������� կ���*�����P��O��8`l��� ����`��ʿϿ��` �	���1p)�H�M� ��phχό���p��x�����V 1��5|�1�!@`y�ŒTHR_INR>0�/�Z"�5d:�MASmSG� Z[�MNF��y�MON_QUEUE ��5�6ӐV~  #tNH�U��qN�ֲ���END�����EXE������BE������OPT�IO������PROGRAM %���%��߰���TA�SK_I,�>�OCFG ά�]���^��DATAu#�����Ӑ2�%B�T� f�x���5��������������,>P�IWNFOu#� ���� ����� '9K]o��� �����/lx�� � ;���ȀK�_�����S&ECNB-�b-&q�&2�/ڝ(G��2�b+ �X,		��=�{���/��@��P4$�0��99)�N'�_EDIT ����W?i?��WERF�L�-ӱ3RGAD�J �F:A�  �5?Ӑ�5Wј6���]!֐��??�  Bz�WӐ<1Ӑn&%�%O�8�;��50!2��7�	�H��l0�,�B=P�0�@�0�M�*�@/�B *�*:�B�O�F�O2��D��A�ЎO�@O	_�,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_�_o �_o�_�_
o�o.o�o jodovo�o�o�o�o�o �o\XB<N� r����4��0� ��&���J������� ����������x� "�t�^�X�j�䟎��� ʟğ֟P���L�6�0� B���f���������(� ү$������>��� z�t��� Ϫ����� �l��h�R�L�^�DX�	���ώ0�� ���t$ :�L��o�
���ߥ��7PREF S��:�0�0
�5?IORITYX�M6}��1MPDSPV��:n" �UT��C�6�ODUCT���F:��NFOG[@_�TG�0��J:?�HI?BIT_DO�8���TOENT 1��F; (!AF�_INE*������!tcp����!ud��8�!�icm'��N?�X�Y�3�F<��1)�� �A�����0� ����������'  ]D�h�������*>��3���9n"OTf�3>�)��2�B�G/�LC���4�;LFJAB,  ���F!/�/%/7/�5�F�Z@�w/�/�/�/�3&�ENHANCE S�2FBAH+d�?�%;�������Ӓ1��1PORT_N�UM+��0����1_CARTRE�@��q�SKSTyA*��SLGS�������C�U�nothing�?�?OO�۶0TEMP �N�"O�E��0_a_seiban|߅OxߕO�O �O�O�O_�O'__K_ 6_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1U@e� v����������Q�<�u�.IVE�RSI	�L��� �disabl�e�.GSAVE ��N�	267_0H771|�h���!�/��9�:� !	^�4�ϐ����e��͟ߟ������9�D�C-Å_y� +1���������ő����Ǻ�URG�E� B��r�WF Ϡ��-��9�W�����l:WRUP_DELAY �=�n�WR_HOT �%��7��/p��R_NORMALO��V�_�����SEMI𓿹�����QSKI%Po��97��xf�=� b�a�sυ�H��ʹ��� ���������&��J� \�n�4�Fߤߒ����� �߲���� �F�X�j� 0��|�������� ���0�B�T��x�f����������ãRBT�IF�5���CVT�MOU�7�5����DCRo���� �T�B׾��C�1bCӏ�&?�q>��ߙ=[H��ٿ��8��^�����ſ*[F��0�KHϘ�� �<
6b<߈�;܍�>u.��>*��<��� �P0���2 DVhz��������,GRDIO�_TYPE  �v��/ED� T_?CFG ��-BH]�EP)�2]��+ �C�u  �/�*��/�?�/%? =�/V?�}?�Ϟ?�� �?�?�?�?�?O
O@O *Gl?qO��8O�O�O�O �O�O�O�O�O_<_^O c_�O�__�_�_�_�_ �_o�_&oH_Mol_o �oo�o�o�o�o�o�o �o"DoIho*j �������. 3�E��f� ���x��� �����ҏ�*�/�N� �b�P���t�����Ο���ޟ�:�+���R'I�NT 2�R��!�1G;� i�{��"x���8f�0 �� ӫ������M� ;�q�W�������˿�� �տ�%��I�7�m� �eϣϑ��ϵ����� ��!��E�3�i�{�a� �ߍ��߱����������A���EFPOS�1 1�!)  x���n#���� ����������/�� S���w����6����� l�������=O�� ��6���V�z � 9�]�� ��Rd��� #/�G/�k//h/�/ </�/`/�/�/??�/ �/?g?R?�?&?�?J? �?n?�?	O�?-O�?QO �?uO�O"O4OnO�O�O �O�O_�O;_�O8_q_ _�_0_�_T_�_�_�_ �_�_7o"o[o�_oo �o>o�o�oto�o�o! �oEW�o>�� �^�����A� �e� ���$�����Z� l�����+�ƏO�� s��p���D�͟h�� ���'�ԟ�o�Z� ��.���R�ۯv�د� ��5�ЯY���}���*� <�v�׿¿����Ϻ��C�޿@�y��e�2 1�q��-�g����� 	��-���Q���N߇� "߫�F���j��ߎߠ� ����M�8�q���0� ��T��������7� ��[�����T����� ��t�����!��W ��{�:�^p ��A�e  �$��Z�~/ �+/���$/�/p/ �/D/�/h/�/�/�/'? �/K?�/o?
?�?.?@? R?�?�?�?O�?5O�? YO�?VO�O*O�ONO�O rO�O�O�O�O�OU_@_ y__�_8_�_\_�_�_ �_o�_?o�_co�_o "o\o�o�o�o|o�o )�o&_�o�� B�fx��%�� I��m����,���Ǐ b�돆����3�Ώ�� �,���x���L�՟p� ������/�ʟS��w������ϓ�3 1� ��H�Z������6�<� Z���~��{���O�ؿ s����� ϻ�Ϳ߿� z�eϞ�9���]��ρ� ��߷�@���d��ψ� #�5�G߁������� *���N���K���� C���g�������� J�5�n�	���-���Q� ��������4��X ��Q���q ���T�x �7�[m� //>/�b/��/!/ �/�/W/�/{/?�/(? �/�/�/!?�?m?�?A? �?e?�?�?�?$O�?HO �?lOO�O+O=OOO�O �O�O_�O2_�OV_�O S_�_'_�_K_�_o_�_ �_�_�_�_Ro=ovoo �o5o�oYo�o�o�o �o<�o`�oY ���y��&�� #�\�������?�ȏ<����4 1�˯u� ����?�*�c�i���"� ��F����|����)� ğM�����F����� ˯f�﯊�����I� �m����,���P�b� t������3�οW�� {��xϱ�L���p��� ��߸������w�b� ��6߿�Z���~���� ��=���a��߅� �2� D�~��������'��� K���H������@��� d�����������G2 k�*�N�� ��1�U� N���n�� /�/Q/�u//�/ 4/�/X/j/|/�/?? ;?�/_?�/�??�?�? T?�?x?O�?%O�?�? �?OOjO�O>O�ObO �O�O�O!_�OE_�Oi_ _�_(_:_L_�_�_�_ o�_/o�_So�_Po�o $o�oHo�olo�oۏ�5 1����o�o�o lW��o�O�s ���2��V��z� �'�9�s�ԏ������ ���@�ۏ=�v���� 5���Y��}�����۟ <�'�`��������C� ��ޯy����&���J� ���	�C�����ȿc� 쿇�ϫ��F��j� ώ�)ϲ�M�_�qϫ� ���0���T���x�� u߮�I���m��ߑ�� �������t�_��3� ��W���{������:� ��^�����/�A�{� ���� ��$��H�� E~�=�a� ����D/h �'�K���
/ �./�R/��/K/ �/�/�/k/�/�/?�/ ?N?�/r??�?1?�? U?g?y?�?O�?8O�? \O�?�OO}O�OQO�O�uO�O�O"_t6 1�%�O�O_�_�_ �_�O�_|_o�_o;o �__o�_�oo�oBoTo fo�o�o%�oI�o mj�>�b� ������i�T� ��(���L�Տp�ҏ� ��/�ʏS��w��$� 6�p�џ��������� =�؟:�s����2��� V�߯z�����د9�$� ]��������@���ۿ v�����#Ͼ�G���� �@ϡό���`��τ� ߨ�
�C���g�ߋ� &߯�J�\�nߨ�	��� -���Q���u��r�� F���j��������� ���q�\���0���T� ��x�����7��[ ��,>x�� ��!�E�B{ �:�^��� ��A/,/e/ /�/$/ �/H/�/�/~/?�/+?��/O?5_GT7 1� R_�/?H?�?�?�?�/ O�?2O�?/OhOO�O 'O�OKO�OoO�O�O�O .__R_�Ov__�_5_ �_�_k_�_�_o�_<o �_�_�_5o�o�o�oUo �oyo�o�o8�o\ �o��?Qc� ��"��F��j�� g���;�ď_�菃�� ����ˏ�f�Q���%� ��I�ҟm�ϟ���,� ǟP��t��!�3�m� ί��򯍯���:�կ 7�p����/���S�ܿ w�����տ6�!�Z��� ~�Ϣ�=ϟ���s��� �� ߻�D������=� �߉���]��߁�
�� �@���d��߈�#�� G�Y�k�����*��� N���r��o���C��� g����������� nY�-�Q�u ��4�X�|<b?t48 1�?) ;u��/;/� _/�\/�/0/�/T/�/ x/?�/�/�/�/[?F? ??�?>?�?b?�?�? �?!O�?EO�?iOOO (ObO�O�O�O�O_�O /_�O,_e_ _�_$_�_ H_�_l_~_�_�_+oo Oo�_soo�o2o�o�o ho�o�o�o9�o�o �o2�~�R�v ���5��Y��}� ���<�N�`������ ���C�ޏg��d��� 8���\�埀�	����� ȟ�c�N���"���F� ϯj�̯���)�įM� �q���0�j�˿�� ￊ�Ϯ�7�ҿ4�m� ϑ�,ϵ�P���tφ� ����3��W���{�� ��:ߜ���p��ߔ�� ��A����� �:��� ��Z���~�����=� ��a���� �����MASK 1����������XN�O  ���� MOTE  �R_CFG �Y�����PL_RA�NGUP���O�WER ���� �A��*SY�STEM*P�V9�.3044 �1�/9/2020 �A � ����RESTART_�T   , �$FLAG� $�DSB_SIGN�AL� $UP�_CND4��R�S232r �� $COMM�ENT $�DEVICEUS�E4PEEC$P�ARITY4OP�BITS4FLOWCONTRO3?TIMEOUe6�CU�M4AUX�T��5INTER�FACsTATUj� KCH� t $O�LD_yC_SW� 'FREEF?ROMSIZ ��ARGET_DI�R 	$UP?DT_MAP"� TSK_ENB"�EXP:*#!jF�AUL EV!�RV_DATA��  $n E��   	$VA�LU�! 	j&G�RP_  � {!A  2� �SCR�	� �$ITP�_�" $NU�M� OUP� �#T�OT_AX��#D�SP�&JOGLI��FINE_PC�d�OND�%$�UM�K5 _M�IR1!4PP TN�?8APL"G0_EXb0<$�!� 814�!{PGw6BRKH��;&NC� IS :�  �2TYP� �2��"P+ Ds�#;0B�SOC�&R N�5DUMMY164�"�SV_CODE_�OP�SFSPD__OVRD�2^�LDB3ORGT-P; LEFF�0<G�� OV5SFTJR3UNWC!SFpF5�%3UFRA�JTO~�LCHDLY7RECOVD'� �WS* �0�E0RO��10_p@  � @��S NVwERT"OFS�@9C� "FWD8A�D<4A�1ENABZ6�0�TR3$1_`1F�DO[6MB_CM��!FPB� BL_MP��!2hRnQ2xCV� "' } �#PBGiW|8AMz3\P��U�B�__M�P�M� �1�AOT$CA� �PD�2�PHBK+!:&a�IO�4 eIDX+bPPAj?a$i�Od7e�U7a�CDVC_DBG"�a;!&�`�B5�e1�j�S�ey3�f�@ATIO� ���AU�c� �S&�AB
0Y.#0 �D��X!� _�:&?SUBCPU%0SIN_RS�T, �1N|�S�T!�1$HW_C1�"]q.`<�v�Q$AT! � ��$UNIT�4|�p�pATTRI= ��r0CYCL3N�ECA�bL3FLT?R_2_FI9a7��c,!LP;CH�K_�SCT>3F�_�wF_�|8��zFqS+�R�rCHAGp��y��R�x�RSD��@'�1E#&7`_T��XPRO�`@S�E�MPER_0�3T�f�]p� f��P�D�IAG;%RAIL�AC�c4rM� LOh�0�A�65�"PS�"b�2 -`�e�SPR�`MS.  �W�Ctazf	�CFUNC�2��RINS_T�.!(�w��� S_� �0�P�� 	d���WARL0bCBL'CUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!2��8�3�TID�S���!� $CE_R�IA !5AFDpPbC~��@��T2 �1C9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@H�RDYOL1	PRG�8�H��>1(�ҥM�ULSE =#Sw3.��$JJJ6BKG�FKFAN_ALMsLV3R�WRNY��HARD�0+&_P� "��2Q���!�5_,�@:&AU�Rk��?TO_SBRvb���� ƺ�pvc�޳MPINF�@�q�)�N��REG'd~0V) x0R�C�1DAL_ �\2FL�u�2$M@Ԑ(�#S��P� `�6g�CMt`NF�qsONIP�q5�IPP� 9a$Y��!�"�!�� �o3EG0P��#@��AR� �c��52�����|5AX�E�'ROB�*REMD�&WR�@�1_=݆�3SY�0ѥ0_�S�i�WRI�@�ƅpST�#��0*@� �q!	���3��� B� �At��3�D�POTO�9� �@ARY�#��0!��d�!1FI�0��$LINK��GkTH�B T_����A��6�"/�XY�Z+"9�7G�OFF��@�.�"���B� l����A3$ ��FI�p���4�4l��$_Jd�"(B�,a������8�"q�������Ck6DUtR��94�TURT�!XZ�N����Xx��P��FL/�@s��l��P��30�"Q +1� K
0M:$�5�3]q7�SuD�Sw#ORQɆ�!�����Q7�
�0O[�ND�=#�!�#�1OVE8��M ���R��R��Q�!P.!P! OAN }q	�R����990�  �brJ9V����Lv�!ER1��	8�!E�@n D�A��p�嘕Ă���v�AX�C�"��`�q� s���0~3� ~F�~e�~�~E�~1��~Ҡ{Ҡ� Ҡ�Ҡ�Ҡ�Ҡ� Ҡ�Ҡ�Ҡ�!)oDEBU}s$x�`��삼!R*�AB��a8A2V`|r 
�"�c���%�Q7� 7�173�7F�7e� 7�7E�����.��LAB����yp��cGRO�p��}��PB_ҁ ��1C���ð�6�1���5���6AND��8p�a3���-G �Q����AH�PH�p2�NTd��Cs@VEL؁�}A��F?�SERVEs@��� $����A!�!�@POR}�KP��b�A �B���	���$�BTRQ�
��CH��@
�G��2	��Eb��_  qlb��Q�ERR��RI�P�@�FQTO	Q�� L�}��YV�ĀG�E%�\ ��CRE�  �,�A�EP
�RA~�Q 2 d�Rr7c�D�A ���$F ׂ��m ��COC��P � 8[COUNT��ђSFZN_CFG�A 4�p%��rT\zs�a�#`pJp�q��&c�� �� MGp+����`�OGp�eFAq����cX8еk�ioQ��'ђ�Dp8�Pz���H�ELA�-b� 5��B_BASN\RSR$�`�2ӑS��L�!p1�W!p2�Dz3Dz4Dz5Dz6�Dz7Dz8�WqROaO���P�1�NL��� �AB�C
�"pAC-K�&IN�PT+�W��U��	�k��y_PUX8�~�|�OU�CP���%�s�Vl���YTPFWD_KARKQL-�:PRE�D�P����QUE$�Ā9 )���~���IU��#s�/���@�/�SEM�1ǆ1�A�aST�Y�tSO����DI��q��Qc��X��_T}M9�MANRQ ��/�END��$K�EYSWITCH�2�G����HE)�BoEATMz�PE��CLEJR���0x�UF��F��G�S�DO_�HOM��Oz��pEFPR��SbJіЊ�uC��O��7P�QO�V_M��}�c�IO#CM���1�Bs;HK�� D,�&�a`U2R��M��a�r �+�FORC*�WA�R䢞�tOM�� � @�$�㰰U���P�1��g���3���4��S�POW�L�z��R%�UNLO��0T�ED�� � �SNP��S�.b 0N�ADD|a`z�$SIZ*��$VA�0�UMULTIP�rj`����Az� � A$��ƒ���SQc�1CFPv�FRIF�r�PSw���ʔf�N=F#�ODBUx�R@�w������F��:�IA`h����������S"p>�� �  �cR�TE���SGL.�T�x�&C`Gõ3<a�/�STMT��`ÙP����BW9 0�S�HOWh�qBANt�TPo���E���h��PV_Gsb; �$PC�0�P�oFBv�P��S�P��A�p���PVD���rb� �+QA002D.ҝ�6�@��6ױ�6׻�6�54�U64�74�84�94�A4�B4و�6ׇ17�}�6�F4� ��@������Z����t�1��1���1��1��1��1���1��1��1��1���23�2@�2M�2�Z�2g�2t�2��2���2��2��2��2���2��2��2��2B��33����M�3Z�U3g�3t�3��3��U3��3��3��3��U3��3��3��3��U43�4@�4M�4Z�U4g�4t�4��4��U4��4��4��4��U4��4��4��4��U53�5@�5M�5Z�U5g�5t�5��5��U5��5��5��5��U5��5��5��5��U63�6@�6M�6Z�U6g�6t�6��6��U6��6��6��6��U6��6��6��6��U73�7@�7M�7Z�U7g�7t�7��7��U7��7��7��7��U7��7��7��7���m�VPv�U�B# �@�09r
�1����A x �0R����  �BM�@RXP�`�4Q_�PR�@P[U�AR��DSMC���E2F_U��=A �SYSL�P>�@ �  �ֲ >g�������iD��VALU>e�pL�Az�HFZAID_L����EHI�JIh�$F�ILE_ ��D�d�$Ǔ�PXCSA�Q� h�0!PE_B�LCKz�.RI�7XD_CPUGY!�GY��Ic�O
TR���R � � PW�`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q�T@J��U�Q�T�Q�UH���T`�T��T2L�_�LIz�  ��pG_OT�P�_EDIU�A�T2�`7c ?bة�pBQ�h����TBC2 �! �%�>��P��a�7aFTτ�d݃TDC�PA�N`�`aM�0�f�a�gTH��"U��d�3�gR�q�9�ERVEЃt݃�t	�.`BC�p�` "X -$EqLENЃRt݃Ep�pcRAv��Y@W_A�tS1Eq�D2�wMO$?Q�S���pI�.B`�A�y�4Ep�{DE�u���LACE �CCqC�.B��_MA�p�v��w�TCV�:��wT,�;�Z�P�Ҡ�s�~��s�J�A�M����J���u)ā�uQq2ѐ����݁�s�JK��V�K������	���J�����JJ�JJ�AAL�<��<��6��:�5�cm�N1�a�m�,��DL�p_�\�Q�ApCF
�#{ `�0GROU�@(J�Բ��N�`C^�Ȑ?REQUIRrÀ�EBUu�Aq��$T�p2"��Bp薋a�	��d$ \?@qhA�PPR��CLB
u$H`N;�CLO}`"K�S�e`��u
�aI�% �3�M�`�l���_MG񱥠C� �"P����&���BR=K��NOLD����RTMO6a�ޭ��	J6`�P>��p��p@��pZ��pc��p6+��7+�<�B� @r�d&�� �lr��x������PATH���������qx�����%0A��SCAub��<�6��INDrUC�p�qZ�C�UM�Y�psP����A q/ʤ��/�E�/�PAYLO�A�J2L�0R_AN�ap�L�Pz�v��jɆ���R_F2LgSHRt��LO{��R�������ACRL_�q�����b�d�9H�@B$H��"�oFLEX>�P�`J�f' P(��o�o�+�p?qJDu( :Qcv�p�����fe��po��|F1 ���-������]�E��*�<�N� `�r�����4�Q����� ��A�c���ɏۏ���	T��2�X:A��� ��������)�;� ?�H�6�Z�c�u�����9>Ѭ�) ��`��0˟ݟ�`�0ATF�𑆢�EL���a��J��(��JE۠CTR��A�TN�1�HAND_VBBq>ѯ@�* $���F2���d�CSW�R�����+� $$M�����0ˡ�@ڡ������A�@ g����A)��A���@
˪A٫A� ��`P�˪D٫D�PȰG�P�)STͧ�!ک�!N�DY�P9���� #%��Fp���Ѫ���i� ���������P3�<�@E�N�W�`�i�r�	�Ҏ�, ��ԓ� �n�5m��1ASYIMص.@�ض+A������_`��	�� �D�&�8�J�\�n�Ju�&��ʧC�I��S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R��&T ��3TWV�͢���&��ߪU��/�7ӂ��03HR`ta-��QLQ�1�DI��O�T8w��P��. ; *"IAA*���$aG�2C�2cJ�$�H��P �/ � �M�E�� Mb�R4AT�PPT�@� ��ua�����P�l@zh�a�iT��@�� $DU�MMY1E�$P�S_D�RF�  t���f3�FLA���YP���b}c$GLB_T��Uuu`�1�=Ѓ�EQa0 XX(���ST�����SBR�PM21_�V��T$SV_E�R��O_@KscsCL�pKrA��O'b�PG�L�@EW��1 4\��a$Y|Z|!W�s怯��AN`�� �sU�u2 ���N�p�@$G�IU}$�q �1� �q�p��3 qL���v^B}$F^B�E�vNEAR��N�K�F8���TANC�K� �JOG���� 4�$�JOINT���� �y��qMSET��5�  �wE�H�� S��u�� ��6�k  MU��?���LOCK_FO�����PBGLVHG�L�TEST_X9M>���EMPt���q�r̀$U�Ќ�r��22���s,�3����Ҁ,�1MqCE����sM� $KAR���M�STPDRA8�pj�a�VEC��{��e�IU,�41�HE�ԀTOOL㠓Vv�RE��IS3��r��6N�A�ACH����5��O�}c�d3ڲ��pSI.� � @$RAIL_�BOXE��ppR�OBO��?�pqHOWWAR*���`�ROLM�bB����S��
�5�0O_�F� !ppHTML5�Q����С2�pڑ��7m�
�R��O��8���v��z�ZЎsOU��9 tpp(�14A��̀��PO֡%PIP��N��
�ڑ�S�,�����CORD�EDҀް̠5�XTL��q)~�� O4` : D pOBP!"Ҁ{�j��cppj�^@$SYSj��ADR#�Pu`TC}H� ; ,��SEN�RZ�Aف_�t�״�>���PV�WVAPa< �� p��r�UPRE�V_RT]1$E�DIT�VSHW�R�7v;���q��@D_`#R�+$HEADoA�Pl��A$�KE�q�`C�PSPD��JMP���L�U
`R��dQ=r�O�϶I�S#�CiNE��$_T�ICK�AM��~���HN-q> �@t������_GP8��[�STYѲ�LOq�r��Ҩ��?�
�Gݵ%$����t=7pS !�$Q��da�e!`�fP�0�SQUd� ��b�ATERCy`�q�p=S�@ �pCp@����d�%Oz`�mcO�IZ�d�q�e�aPRM��a8����sPUQH�_DO=��ְXS��K�VAXiIg�f�1�UR� ���$#�Е��� _,����ET��Pۂ�� �5`o��6g�A�!�1��d9�2;� �SR|Al �о���#��5�� #��#�)#�)i�>' i�N'i�^&{����){�H���2��C����C���WOiO{O�D��SSC�p B hppD1S(�k��`SP`�ATL �I����~�bADDRES��=B'�SHIF��"��_2CH#��I\&p��TU&pI�� C͢CUST�O��~�V��IbD�Ȳ,��0
�
ⶲV�X�R`E \�����f�7��tC�#	���F��irt��TXSCREE�l�F�P��TIN!A�s�p��t������0G T��fp,� ��eqBp&uᦲu�$#�RRO'0R���}��!��HaUE��H ���0���`S�q��RSM�k�UV����V~!�PS_�s�&C�!�)�'C��Cǂz"�o 2G�PUE�4�Ibvr�&8�GMT
jPLDQ��Rp�z�/BBL_�W�`R`�J �f�>2O�qJ2LE�U3"�T4�RIGH^3BRD<xt�CKGR�`�5�TW��7�1WIDT�H�H����a�a��o�UIu�EY��QaK d�p��A�J�z
�4�BACKH�h�b�5|qX`FOD�nGLABS�?(X`yI�˂$UR(��9@���0^`H4! 'L 8�QR�_k��\B_`R�p͂����a��IAO�R`M�$�w0Uj0�CRۂM��LUM�C��� ER�V��p�0P<��4NV`��GE=B#���L]�t�LP�E��E��Z)Wj'Xz'XԐ�&Y5$[6$[7$[8 	R���3�<���fԑ�ŁS��M�1U{SR�tO <��b^`U�r�rFO
.�rPRI��m�����PTRIP�m��UNDO��P�p��`m�4���#���� QWB�P7�G s�Tf�H�&RbOS�agfR��:">c��.qR��s�~�b$*�<eUQ.qS�o�op�#R)�>cOFF����pT� �cOp G1R�t/tS�GU��P.q��JsE�Tw�1SUB*� �f�E_EXE��V���>cWO>� U2�`^g��WA'��P�q!@� V_DaB�s�pJ�>`RT�`�
�V�Q�r��OR���uRAU��tT��ͷ�q_���W 9|%�͸OWNA`޴$SRCE � ���D��\��MPFI8A�`��ESPD�� ����C���Gƒ�r-�5��!X `�`�r޴���COP�a	$��C`_w������rCT�3�q���q�ƒ�0��@� Y~"SHADOW�����@�_UNSCAp��@��4M�DGDߑ��EGAC�,���PPG�Z (�0NO�@�D<�PE��B��VW�S�G|���![ � ���VEE#�aڒANG��$��c薴cڒLIM_X�c��c� � ���#��`� ��b�VF� �s�VCC�jв�\ՒC{�RA�lצ���RpNFA���%�E��Z2`G� ^0[�C`�DEĒ��� STE Q1���@�ꁻ@I��`�+0����`����P_A6�r���K��!]� 1Ҡ���A��\��сCPC�@�]�DRIܐ\�͑V�#Ѐ���D�TMY_UBY�T���c��F!���Y��$����P_V�y��LN�B�MQ1$��DEY���EX�e��MUj��X�M� US�!���P_R��b�P� zߖG��PACIr� ʐf�ᔟ��c�´c��#�EqB��a.28B����^ ܀�GΐP����`C�R~``�_�0�@3!�1zri	�e�R�SW�� p�00��S�6�O�Q�1�A� X�#�E�UEd��00pC�HKJ�`�@p���U� �EAN�ٖp�pXռ�`C�MRCV�!a� ��@O��M�pC«	��s����REF*7
��������/� �P��@���@��b�����_Y��ژ��ۣ�� Q$3����Ӷ�C��$b ����%���Q~��$GROU�  �c�����ʠ]��I�2^0��U` 0�_�I,�o � UL�ա`��C&�rAaB�?�NT����$��� �A���Q��K�L����@õ��A���Q��T na$c t�`MD�p�8�HU���SA.�CMPE F  _�Rr�p@����XS	qVGF|/�b#d, &�@qM�P^0۰UF_C 0!���z �ROh0"�+���@���0C�UR1EB���RI��
IN�p�����d���d��ca�INE�H�y��0V�a-�걗�3�W�������C��i�LO�}�z�p@0�!�QNSI���݁���c$&�c$&.�X�_PE-YW+Z_IM�ڒW�I�$��" �+R�'rRSLNre �/�M
`R�RE�C7�Gd� ۰�̵ҭ�q����u ��Ȑ������S�_P�VnP m�V�IA�vf �~pHkDR�p�pJO�P���$Z_U�P��a_LOW��5�1J�dA��LINubEP?�tc_i�1�1���@�G1@�V��xg 5X�P�ATHP X�CACH$�]E��yI��A��{�C)�ID3F�A�ETD�H��$H�O�pO�b@�{��d6�F�����p�PA3GE�䁀VP�°��(R_SIZ��2TZ�3�-X�0U�q�MP\RZ��IMG���sAD�Y�MRE���R7WGP��8�p��ASYNBUF�VRTD�U�T7Q�LE_2D-��U�J�`CҡU1��Qu���UECCU��VE�M��]EDb�GVIR�C�Q�U�S�B�Q�L�A��p�NFOUN^_�DIAG�YRE�GXYZ�cE�W� �h8�dpqa`T��2IM�a�V|be��EG/RABB��Y�aЗLERj�C4���FC-A�6504x��7u�$�@G��h��`�CKLAS_@l�BA��NN@i  G��T��� @ݲմ$BAƠwj �!q�eb��u�TYSp�H����2��I��t:b�f��B)�EVE����PK���fx6��GI�pNO��2����#�HO����k � ���
8�Pbi�S�0ޗ��ROⓟACCEL?0=���VR_�U7@�`���2�p��AR��PA蹀̎K�D��REM�_But *�#�J�MX �l�t�$SSC�U���!#����QN@m � �S�P�NS��LEX�vn T�ENA�B 2�W@��FLDRߨFI�P�t�ߨ�(Ğ��2P2HFoO� ��V
>Q MV_PI��@8T@󐉰�F@�Z�+�#��8��8#��GAB���LsOO��JCBx���w"SCON(P�P�LANۀ�Dp�3F �d�v�9PէM��Q ;����SM0E�ɥ� 8ɥWb72$`<�8T���,`RKh"ǁV�ANC��@AR_Ou N@p (�-#<#@c��c2� w�A/�N@q 4������`p	�^���r hn�p��1^�&OFF`�|�p�`��`�DEA��
�P,`SK�DM�P6VIE��2q �w��@���rs <C {���4���r�{7��D���}qC�UST�U��t� $G�TIT1�$PR\��OPyTap ��VSF��
�su�p�0`r&�]��SMOwvI�d|�ĄJ�����eQI_WB��wI���� x@O3�@�XVRx�xmr��T�� ��ZABC��y� op����)�
	���ZD$�CSCH��z Lu����`�2��%PC ��7PGN� ��<��A��_FU�NH��@ �Z�IPw{I��L�V,SL��~�  �ZMPCF���|��E����X�DM�Y_LNH�=���M�|��} $x�A� ]�CMCM� EC,SC&!��P��? $J���DQ������������±�_�Q,2����UX|�a\�UXEUL� �a������(�:�(�<J���FTFL��w�n�Z�~?@L+�6� f���Y@�Dp  8 �$R�PU��> EgIGH����?(��iֱ��0��et� a�a�����$B�0��0@�	�_SHIYFD3-�RVV`F�@&��	$5��C�0��@&!������b
�s4x�uD�TR��9V����SPH���!�� ,������� ��4A�RYP���%�����%���"P�%!���H�(UN0���"�2������K��q0G�SPDak�� ��P��O����0X��Я�"!�NGVER`q �iw+I_�AIRPURGE�  i  �i/�F`E�Tb� ΋+  � h2IS_OLC  �,�"�!���!�%��P+Y�_/*OB��Dm��?@�!H771  34 n?�?�9� `�E/#�)�x� S232�� �1i� L�TEk@ PEN�DA�341 1D�3<*? �Maintena�nce Cons� B�? F"O,D?No UseMJO OnO�O�O�O�O2�2GNPO;/" 19%��1CH=� ��-Q		9Q_!�UD1:___RSMAVAIL/��/%�A!SR  �+��H�_�P1�oTVAL.&����P(.�YVL�}� 2�i�� D��P 	�/_oUQNo �orci�o�g�o�o�o �o�o*,>t b������� ��:�(�^�L���p� ������܏ʏ ��$� �H�6�X�~�l����� Ɵ���؟�����D� 2�h�V���z������� �ԯ
���.��R�@� b�d�v�����п���� ���(�N�<�r�i��$SAF_DO_PULS. jQp����CA� �/%��&0SCR ��`}X��0�0
	14�1IAIE��@�0 vo$�6�H� Z�l�~�ߢߴ�����X�����HS��2%�����d1�(�8�qrb��� @�"@k�}���T�h� J`����_ @��T7 �����#�0�?T D��0�Y� k�}������������� ��1CUgyx�O�Ef������  �5;G�o�� 1p�U��
�t��D�i�������
  � ��*������g y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O<A���`OrO�O�O�O �O�O�O�O?O�_._ @_R_d_v_�_�_�_�_�Q _�R0MJT o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏJO��'�9�K�]� o�������_ɟ۟� ���#�5�G�Y��_�U �_�ҙ�����ϯ�� ��)�;�M�_�m��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0�B�T�f�;�?�q� ������������,� >�P�b�t������������������Y��	�12345678�1h!B!S����F��� ��������������  ��;M_q� ������ %7I[l*�� �����//1/ C/U/g/y/�/�/�/n ��/�/	??-???Q? c?u?�?�?�?�?�?�? �?O�/)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_O_�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o p_�o�o�o/A Sew����� ����o+�=�O�a� s���������͏ߏ� ��'�9�K�]���� ������ɟ۟���� #�5�G�Y�k�}�����D����s�կ�w����0�L�CH � Bpw�   ��=�2�� _} =�
��?�  	�o�ί ��ǿٿ���r������@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖ�%Ϻ� ��������&�8�J� \�n���������@�����"�Q�*�����;�<M���D���?  �]�w��*�Z򛱛�t  �d�����*�`*���$SCR_GRP� 1*P�3� � ��*� 6�	 �
��<�+*��'UC|@��,y�yD� W�!��y�	M-1�0iA/7L 1�23456789�0��� 8��cMT� � �
�	dL��	Č� N
���Y���y"�
M_	P����� ,�G�H�
 ��� 1/@A/g/y/H�ߙ!T/�/P/�/3��+��.�/B�S��,?*2�C4&Ad�R?  @0s�j5N?�7?��7&2�R��?}:&F@ F�`�2�?�/�?�? OO-OSO>OwObO�O =j1�2�O�O�O�O�DB��O�O;_&___J_ �_n_�_�_�_�_�_o �_%o�5j�eSgxo6���uo�o�b�1�B�|3�oh0�4j9j9B� w�$Y̯@HtA�Nhcu�/��%pp�drsq  ����z�q�x�\ �� (&�*� 2�D�V�oz�e��������ECLVL  �����iqpQ�@��L_DEFA�ULT ���s�փHOOTSTR�qq���MIPOWERF���H���WFD�O� �RV?ENT 1ɁɁ�� L!DU�M_EIP������j!AF_IN�E‧���!FT$}�֞����!-/�� ��F�!RPC_MAING��)��5���Y�VIS�b�t����ޯ!TMPѠPUկ��dͯ�*�!
PMON_�PROXY+���e �v��D���fe�¿�!RDM_SR�Vÿ��g���!�R,*ϑ�h��Z�!%
[�M����iIϦ��!RLSYNÇ���8����!gROS|���4���>�!
CE�MT'COM?ߓ�k-ߊ�{!	S�CONS�߲��ly���!S�WOASRCݿ��m��v"�!S�USB#��n�n�!STMC��o]��� ��ѳ����,���P��V�ICE_KL �?%d� (%SVCPRG1S�����2�������o��"��4������5"��6;@��7ch������9�� ��%�������� 0����X����� -���U���}� �� /���H/��� p/���/��F�/�� n�/��?��8? ���`?��/�?��6/ �?��^/�?��/X�j� ��q���#OhO��lO�O {O�O�O�O�O�O�O _ 2__V_A_z_e_�_�_ �_�_�_�_�_oo@o +odoOo�o�o�o�o�o �o�o�o*<` K�o����� ��&��J�5�n�Y����}���ȏ���^�_�DEV d���MC:�4����GRP 2�d���bx 	� 
 ,V���s�Z����� �������ߟ�� @�'�9�v�]��������Я����۫Y��"��ܯ�1�4� ]���j�����˿Ӵ� ������0��T�;� Mϊ�qϮ��[�!��� ���ߡ�K�!�^�p� ���s�Y��ߩ����� 
���@�'�d�v��y��^�������� ��%��I�0�Y��f� ��������������� 3��T7]�e� ���z����� 1Ag"�r�@��=����� �!/G/���R/�/�/ �/�/�/"�/�/?? C?*?<?y?`?�/�f? �?�?�?�?�?-OOQO 8OaO�OnO�O�O�O�O �O_�O)_;_"___�? �_�_L_�_�_�_�_�_ o�_7oo0omoTo�o xo�o�o�o�o�o! x_E�oU{b�� ������/�� S�:�w�^�p�����я��d �X�ZI�6 r 	 �@Z��0�+�A����d�BjBA�=��������B����AZ.�A����+�A.��Q�B�����5\��i6�A��u��'��ǎ%�Ꮛ�%�PEGA_BAR�RA_ESTEI�RA����X�T����?=��=�X��7
�?��>�A����?������&����������AxP��f���U�'A�j���´�B��:�<�3�����jB]+a��T��%�T�腯d�ʐ���>�p�c?��7�Գ�T@6��A�_���0n�����·�Ak���۸I�K9�FA�G�����B!v,�-���C3�����pBM�>�#�b��(�Y�������HX��?L!���Q��B���AJߤ�Xk�@f�D3��O�A���������Yw���.B��B�;��C�H�z�B�?���6���-Ϙ������n��=]����V@����?,����Ö� վ���eAk�������OY�A��ㇾ��AB��J�;%�C$�4�aƿBXZ�9���
���ߘ��~��� �ԭ(��?^_��-\¯ԡ���گ���+������������ߔ�mᢧ��*נ�6�C>�ԯb���z���
��BM����s��x�U<~�߯7@6|=��C��$�6��� N�@���b�G���L��}������x7���~K@����V�+A>r�rF���������Y@+�@��<B��|�A��F����B)���,o�?ɇ���~0��0~�6�Z� Q������������Aߍ�]ܖ�A����ܺ����2[�����>�ȥA���=�³�NB ��$�w?�d�j��to�7\��
�.�%��Z�����A������*�@Ve��B� ������YN�#���BD�	����9A����gB#
q��3��C4#���,?[BVM����COLO�CA_PRENS|���X�\{B*3Vhz��������/
&�M�@/(/:/L/^/p&�z/��/�/�/�/�/X�N�&v��*�@�n�4B-N���vB��������9���z��@�k'@л���آjA���̶�QB!dD���R?�o��^��CU�@Z??O~?�?uO{B� O�O�O�O�O�O�O  _G__x_f_�_ �_�_�_�_&_L_o\_ �_Po>otobo�o�o�o �_�o"o�o�o&L :p^��o��o� ��� �"�H�6�l� ����\�Ə���؏ ����D���k���4� �������ԟ
�L� 1�C������d����� �����$�	�H�ү<� *�L�N�`��������� � �����8�&�H� J�\ϒ�Կ�������� �����4�"�Dߚ��� ����j��߲������ ��0�r�W�� ��� ����������J�/� n���b�P���t����� ����"�F���:( ^L�p����� � 6$ZH ~���n�j� /�2/ /V/�}/� F/�/�/�/�/�/
?�/ .?p/U?�/?�?v?�? �?�?�?�?OH?-Ol? �?`ONO�OrO�O�O�O O4O_DO�O8_&_\_ J_�_n_�_�O�_
_�_ �_�_o4o"oXoFo|o �_�o�_lo�o�o�o�o 
0T�o{�oD �������,� nS�����t����� Ώ���4��+��� ޏL���p�����ʟ� �0���$��4�6�H� ~�l����ɯ����� � ��0�2�D�z��� ���j�Կ¿���� 
�,ς���yϸ�RϬ� ���Ͼ������Z�?� ~��r�߂ߨߖ��� ����2��V���J�8� n�\�~�����
��� .��"��F�4�j�X� z�������������� B0f���� VxR��� >�e�.��� ����/X=/| /p/^/�/�/�/�/�/ �/0/?T/�/H?6?l? Z?�?~?�?�/?�?,? �? OODO2OhOVO�O �?�O�?|O�OxO�O_ 
_@_._d_�O�_�OT_ �_�_�_�_�_oo<o ~_co�_,o�o�o�o�o �o�o�oVo;zo n\����� �����4�j�X� ��|����ُ���� ����0�f�T���̏ ����z��ҟ���� �,�b�����ȟR��� ���ί���j��� a���:���������ܿ ʿ �B�'�f��Z�� jϐ�~ϴϢ������ >���2� �V�D�fߌ� z߰�����ߠ�
��� .��R�@�b���߯� ��x��������*�� N���u���>�`�:��� ������&h�M�� �n����� �@%d�XF| j�����< �0//T/B/x/f/�/ �/�//�/?�/,? ?P?>?t?�/�?�/d? �?`?�?O�?(OOLO �?sO�?<O�O�O�O�O �O _�O$_fOK_�O_ ~_l_�_�_�_�_�_�_ >_#ob_�_VoDozoho �o�o�oo�o�o�o�o �oR@vd��o � ������ N�<�r�����b�̏ ����ޏ ���J��� q���:�����ȟ��� ڟ��R�x�I���"�|� j�����į���*�� N�دB�ԯR�x�f��� ������&����� >�,�N�t�bϘ�ڿ�� ����������:�(� J�p߲ϗ���`��߸� ����� �6�x�]�o� &�H�"��������� �P�5�t���h�V�x� z���������(�L� ��@.dRtv� � �$�< *`Np���� ���//8/&/\/ ��/�L/�/H/�/�/ �/?�/4?v/[?�/$? �?|?�?�?�?�?�?O N?3Or?�?fOTO�OxO �O�O�O�O&O_JO�O >_,_b_P_�_t_�_�O �_�_�_�_�_o:o(o ^oLo�o�_�o�_ro�o �o�o�o 6$Z�o ��oJ����� ��2�tY��"��� z�����ԏ�:�`� 1�p�
�d�R���v��� ��П���6���*��� :�`�N���r����ϯ �����&��6�\��J���¯������$SERV_MA_IL  �����ʴOUTPU}Tո�}@ʴRV 2j�;  � (r�������=�ʴSA�VE���TOP1�0 2� d? 6 rƱ�� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b�0t�����n�YPY���FZN_CFG ;f��=���J���GRP 2���g� ,B �  A �D;�� B �  B�4=�RB21�I�HELL�� f�e�)�*�=����>�%RSR�� ����&J 5G�k�������.�  ��/>/P/"\/1�1X/1�2��U'&"�2�dh,g-�"EH�K 1S  �/�/�/�/#?L?G?Y? k?�?�?�?�?�?�?�?��?$OO1OCO?OM�M S�ODFTOV_ENBմ��e��"OW_RE�G_UI�O�IM�IOFWDL~@x�N�BWAIT�BA�)��V��F��YTIM�E���G_VA԰_�A_U�NIT�C~Ve�LC��@TRY�Ge��ʰMON_ALI_AS ?e�I%�he��oo&o8oFj �_io{o�o�oJo�o�o �o�o�o/ASe w"������ ��+�=��N�s��� ����T�͏ߏ��� ��9�K�]�o���,��� ��ɟ۟ퟘ��#�5� G��k�}�������^� ׯ�����ʯC�U� g�y���6�����ӿ� �����-�?�Q���u� �ϙϫϽ�h������ �)���M�_�q߃ߕ� @߹������ߚ��%� 7�I�[������ ��r������!�3��� W�i�{���8������� ������/ASe �����|� +=�as� �B����/� '/9/K/]/o//�/�/ �/�/�/�/�/?#?5? �/F?k?}?�?�?L?�? �?�?�?O�?1OCOUO gOyO$O�O�O�O�O�O �O	__-_?_�Oc_u_ �_�_�_V_�_�_�_o�oc�$SMON�_DEFPROG &���Aa� &*SYSTEM*o~bg $JO0d�RECALL ?�}Ai ( �}�=copy md�:pickup_�barra_es�teira.tp� virt:\t�emp\=>10�.109.3.6?2:8460bo�o��o	x};�o�`torno�o�m�oj|zz4vlace1�C�aR��� }}:usumir+ ��h�j�|��w�cprens�oH�������6|��Ï�a�ԏe�w�
�<�furad��<��o������v%�sem_recep1���ʟZ�0l�~����fco-�?�pQ����� }9u�drop*�defeit5�ɮׯh�z�2�7�.�_15�ɏ`W��������_2���ſ׿h�z���_3�3�E�W������x�yzrate 61�� ����]�o߁�:��
�11 C�:� L�������&߸����[�m���frs:�orderfil�.dat��mpbackA�V�W�������-tb:*.*���ʭ��\�n����1x��:\&���8�S�PT�������2��a�����ԣ��as���61 (:L����ϣ12624 ��^p�� ��5G���!�84:15972���]/o/�/��tpdisc 0'/2 9/K/�/�/ ?��tpconn 0�ذ/�/�/e?w?
? �â�+�,,U?�?�?�.��?0(�?]OoO�O &�2&PO�O�O_q3�O+-�Ob_t_ �_�?�?4OOO�_�_o O�_;O�_^opo�o�O &o:_�O�o�o _%_ �oI_Zl~�_�_,o �_���o!o�Eo �h�z��o�o2�oU� �����Aӏd� v�����6�Q���� ����=�ϟ`�r������$SNPX_�ASG 2�������3 T��%���Я�  ?���PAR�AM ��^�� �	��PӤ���Ө$�������OFT_KB_CFG  ӣ�����OPIN_S_IM  ����}���������RV�NORDY_DO�  )�U���QSTP_DSBi���ϐ�SR }�� � &#��D�O�O�:�TOP_ON_ERRʿ���o�PTN z�����A���RING_PRM�y�ܲVCNT_GOP 2��!���x 	���ϗ���#���Gߔ�VD��RP' 1��"�8Ѩ� *߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�}�z����� ����������
C @Rdv���� ��	*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?[?X?j?|?�? �?�?�?�?�?�?!OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLoso po�o�o�o�o�o�o�o  96HZl~ ��������� �2�D�V�`�PRG�_COUNTJ�9��{�ENB��}��M��L���_UPD� 1'�T  
k������"�K�F� X�j���������۟֟ ���#��0�B�k�f� x���������ү���� ��C�>�P�b����� ����ӿο���� (�:�c�^�pςϫϦ� �������� ��;�6� H�Z߃�~ߐߢ����� ������ �2�[�V� h�z���������� ��
�3�.�@�R�{�v� ������������ *SN`r����t�_INFO {1�Ҁ� 	 ��3�@�1�?�|��?��9 B���ƓA��&���ߌ��I�@L>�>�` AoB �@{w ?�� �>�@��a� A  %Cj���D���3����7�lB�� ���YSDOEBUG����� �dՉ�SP_PA�SS��B?+L_OG ���� �  a� � �с�UD�1:\;$�<"_M�PCA-셽/�/��x!�/ 쁝&SAV D)��%d!|"��%�(SV�+T�EM_TIME �1D'�� 0Xh������()���#-M7MEMBK'  �сd d/x�?�?�<X|Ҁg� @�?C�O :OJLOmOzI�J
! %@p1�O�O�O �O"3 __$_6_H_Z_l_ �n_�_�_�_�_@�_�_�_o"o\�e1o Vohozo�o�o�o�o�o �o�o
.@Rd`v���O5SK�0��8���?���F�ҀB�H2OJ�}AJ� �`�аA\O����(�O"��Oяb�ݏw_�O? 3 � ��0'#Z� l�~�����Q��Ο������$�C�7o g�y���������ӯ� ��	��-�?�Q�c�u�����������T1SVGUNSPD%%� '%��2M�ODE_LIM #a9"ܴ2�	�� D-۵ASK_?OPTION �9�!F�_DI ENB  U�%f��BC2_GRP 2!�u#o2��N���C���ԼBCCF�G #��*< #6���q�*�N� 9�r�]ߖߨߓ��߷� �������8�#�5�n� Y��}��������� ���4��X�C�|���  t���u����� c���	B-f�. ��4[ ����� �� 02Dz h������� /
/@/./d/R/�/v/ �/�/�/�/�(���/? &?8?J?�/n?\?~?�? �?�?�?�?�?O�?4O "OXOFOhOjO|O�O�O �O�O�O�O__._T_ B_x_f_�_�_�_�_�_ �_�_oo>o�/Voho �o�o�o(o�o�o�o �o(:Lp^� ������� � 6�$�Z�H�~�l����� ��؏Ə��� ��0� 2�D�z�h���To��ȟ ���
���.��>�d� R�������z�Я���� ���(�*�<�r�`� ��������޿̿�� �8�&�\�Jπ�nϐ� �Ϥ������ϴ��(� F�X�j��ώ�|ߞ��� ���������0��T� B�x�f�������� ������>�,�N�t� b��������������� ��:(^�v� ���H���$ HZl:�~� ������2/ / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?P? R?d?�?�?�?t�?�? OO*O�?NO<O^O�O rO�O�O�O�O�O�O_ _8_&_H_J_\_�_�_ �_�_�_�_�_�_o4o "oXoFo|ojo�o�o�o �o�o�o�o�?6H fx���������v&��$TB�CSG_GRP �2$�u��  �&� 
 ?�  Q�c�M� ��q��������ˏ���*�1�&8�d�, �F�?&�	 �HCA�����b��CS�B�I�����V�>���ͪ�n�Ќ�ԝB���333��Bl"t������AÐ��fff:��.�C�����l�?�� ��G�w�R���A&��̧�����@��I�� -���
�X�u�@�R���轿̻�����	V�3.00I�	mt7���*� �%���ֶY��@f�f&� &�H�� �N� �O�  ������ ϏϘ�*�J2�1�'8��Ϥ�CFoG )�uB�Y E������d�9��#��#�I� W��pW�}�hߡߌ��� ���������
�C�.� g�R��v������ ��	���-��Q�<�u� `�r����������� I�cp"4��gR w������	 -?�cN�r ��&������ /</*/`/N/�/r/�/ �/�/�/�/?�/&?? J?8?Z?\?n?�?�?�? �?�?�?O�? OFO4O jOXO�O�O`�O�OtO �O_�O0__T_B_x_ f_�_�_�_�_�_�_�_ �_,ooPoboto�o@o �o�o�o�o�o�o�o( L:p^��� ����� �6�$� F�H�Z���~�����؏ Ə����2��OJ�\� n������������ ��
�@�R�d�v�4� ��������ί���� ү(�N�<�r�`����� ����ʿ̿޿��8� &�\�Jπ�nϐ϶Ϥ� ��������"��2�4� F�|�jߠߎ����߀� �� �߼�B�0�f�T� ��x��������� ���>�,�b�P����� ����v������� :(^L�p�� ��� �$H 6lZ|���� ��/�/ /2/h/ �߀/�/�/N/�/�/�/ 
?�/.??R?@?v?�? �?�?j?�?�?�?�?O *O<ONOOO�OrO�O �O�O�O�O�O _&__ J_8_n_\_�_�_�_�_ �_�_�_o�_4o"oXo Foho�o|o�o�o�o�o �o�/$6�/�ox f������� �,�>���t�b��� ����Ώ��򏬏�� &�(�:�p�^������� ��ܟʟ�� �6�$� Z�H�~�l�������د Ư��� ��D�2�T� z�h���Jȿڿ�� ����
�@�.�d�Rψ� vϬϾ����Ϡ���� ��*�`�r߄ߖ�P� �ߨ���������� &�\�J��n����� ��������"��F�4� j�X�z�|��������� ����0B�Zl ~(������ �,Pbt�D�������  9 # &0/�"�$TBJOP_GRP 2*���  �?�&	H"O#,vV,���� ן� =k% � Ȫ � �� ��$ @ g"	� �CA��&�?�SC��_%g!��"G��"k���/�+=�C�S�?��?��&0%0CR  B4��'??J7�/�/?33�3�2Y&0}?�:;���v 2�1�0-1*�20�6?�?20��7C�  D�!�,� �BL��OK:��Z�Bl  @pzB@�� s33C�1y �?gO  A�zG�2jG�&)A)E�O�J�;��|A?�f�f@U@�1C�Z0z8jO�Oz@���U�O��$fff0R)_;^;7xCsQ?ٶ4)@ �O�_tF�X_J\EU�_��V:�t-�Q(B� *@�Ooh�&-h$oZG Lo6oDoro�o~o8o�o �o�o�o3�oR@lVd��V4�&�`�q�%	V3.{00m#mt7A@��s*�l$!�'�� E��qE����E�]\E���HFP=F��{F*HfF@�D�FW�3Fp�?F�MF����F�MF���F�şF���F�=F����G�G�.8�CW�RD�3l)D��E�"��Ex�
E���E�,)F�dRFBFHF�n� F��F���MF�ɽF��,
GlG�g!G)�G�=��GS5�G�iĈ;��
;W�o�|& : E@Xz&/��&�"�?�0�&=;-E�STPARS  �(a E#HRw�A�BLE 1-V)� @�#R�7� (� �R�R�R�'T#!R�	R�
R�R�T��!R�R�R����RDI��`!���ԟ���
�r�O z���������̯ޮ��	Sx�^# <�����ÿ տ�����/�A�S� e�wωϛϭϿ����� ��;-w�{�_"��6�� 1�C�U���%�7�I��[����NUM  ��`!� �$  ��m���_CF�G .���!@�H IMEBF_T�T}���^#��G�VE�10m�H�]�G�R {1/�� 8��" �� �A�  ������������  �2�D�V�h�z����� ��������/
e @Rhv���� ���*<N `r������ '///]/8/J/`/n/@�/�/�/�/r���_���t�@~�t�MI_�CHANS� ~� ~!3DBGLVLS��~�s�$0ETHE�RAD ?��
w0�"��/�/�?�?�l�$0ROUTq��!�!�4�?�<SNMASKl8~�}1255.2E�s0O�BOTO�st�OOLO_FS_DI}��%�V9ORQCTRL� 0���#��MT �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo&l�OIo8omoq��PE_DETAI�J8�JPGL_CONFIG 6��ᄀ/cel�l/$CID$/grp1qo�o�o/壀�?Zl~ ���C����  �2��V�h�z����� ��?�Q����
��.� @�Ϗd�v��������� M������*�<�˟ ݟr���������̯@�}a���&�8�J�\���^o��c��`���˿ ݿ���Z�7�I�[� m�ϑ� ϵ������� ���!߰�E�W�i�{� �ߟ�.���������� ��A�S�e�w��� ��<���������+� ��O�a�s�������8� ������'9�� ]o����F� ��#5�Yk�}�����`��User Vi�ew �i}}12�34567890 �//,/>/P/X$� ,�cx/���2�U �/�/�/�/??s/�/�3�/b?t?�?�?�?�??�?�.4Q?O(O�:OLO^OpO�?�O�.5 O�O�O�O __$_�OE_�.6�O~_�_�_�_ �_�_7_�_�.7m_2o DoVohozo�o�_�o�.8!o�o�o
.@��oagr lCamera� �o����� �ޢE�*�<�N��h�z�`�������I  �v �)��$�6�H�Z�l� ���������؟���� �2�Y��vP9ɟ ~�������Ưد��� � �k�D�V�h�z��� ��E�W�I5�����  �2�D��h�zό�׿ ����������
߱�W� ދ��X�j�|ߎߠ߲� Y�������E��0�B� T�f�x�߁ulY��� ������
����@�R� d�������������� ��W� iy�.@Rd v�/����� *<N��W��i �������� /*/</�`/r/�/�/�/�/as9F/�/? ?1?C?U?�f?�?�? D/�?�?�?�?	OO-O
�j	�u0�?hOzO�O �O�O�Oi?�O�O
_�? ._@_R_d_v_�_/OAO �p�{,_�_�_oo)o ;o�O_oqo�o�_�o�o �o�o�o�_�u���o M_q���No� ��:�%�7�I�[� m�NEa����ˏݏ ����7�I�[��� �������ǟٟ���� ͻp�%�7�I�[�m�� &�����ǯ����� !�3�E�쟒�9�ܯ�� ����ǿٿ뿒��!� 3�~�W�i�{ύϟϱ� X�����H����!�3� E�W���{ߍߟ����������������  ��L�^�p���������� ��   "�*�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</�N/`/r/�/�  
���(  �@�( 	 �/�/�/�/ �/? ?6?$?F?H?Z?@�?~?�?�?�?�*2� �l�O/OAO�� eOwO�O�O�O�O��O �O�O_TO1_C_U_g_ y_�_�O�_�_�__�_ 	oo-o?oQo�_uo�o �o�_�o�o�o�o ^opoM_q�o�� ����6�%�7� ~[�m��������� ُ���D�!�3�E�W� i�{�ԏ��ß՟� ����/�A�S���w� ����⟿�ѯ���� �`�=�O�a������� ����Ϳ߿&�8��'� 9π�]�oρϓϥϷ� ��������F�#�5�G� Y�k�}��ϡ߳���� ������1�C�ߜ� y������������� 	��b�?�Q�c���� ����������(� )p�M_q������0@ �������� ��#�frh:\tpg�l\robots�\m10ia4_?7l.xml�X j|�������.��/1/C/U/ g/y/�/�/�/�/�/�/ �//?-???Q?c?u? �?�?�?�?�?�?�?
? O)O;OMO_OqO�O�O �O�O�O�O�OO _%_ 7_I_[_m__�_�_�_ �_�_�__�_!o3oEo Woio{o�o�o�o�o�o �o�_�o/ASe w�������o ��+�=�O�a�s����������͏ߏ��I �<<w  ?�� 4��,�N�|�b����� ��ʟ�Ο���0�� 8�f�L�~���������������(�$T�PGL_OUTP�UT 9����;� $�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ�����$�����2345678901��� � 2�D�V�^����υߗ� �߻�����w����'�9�K�]���}g��� ������o����1� C�U�g���u������� ����}���-?Q c������� ��);M_q 	������ �%/7/I/[/m/// �/�/�/�/�/�/�/? 3?E?W?i?{??%?�? �?�?�?�?O�?OAO SOeOwO�O!O�O�O�O��O�O_�O� $$Ӣ��OW=_o_ a_�_�_�_�_�_�_�_ �_#ooGo9oko]o�o �o�o�o�o�o�o�oC5g}��� �����}@���"�� ( 	 iW�E�{�i����� Ï��ӏՏ���A� /�e�S���w������� �џ���+��;�=��O���s����Ƹ  <<\ޯ� )�ͯ�)��M�_��� ʯ����<���ؿ��Ŀ � �~�$�V��Bό� ��x�����2ϼ�
ߤ� ��@�R�,�v߈���p� ����j�������<� �߬�r������ �����`�&�8���$� n�H�Z���������� ����"4Xj�� R��L���� |Tf �� v��0B//� &/P/*/</�/�/��/ �/h/�/??�/:?L? �/4?�??n?�?�?�? �? O^?�?6OHO�?lO ~OXO�O�OO$O�O�O �O_2___h_z_�O �_�_J_�_�_�_�_o�.o��)WGL1�.XML�cm�$�TPOFF_LI�M Š�p��{�qfN_SVy`�  �t�jP_�MON :����d�p�p2miS�TRTCHK �;���f~tbVT?COMPAT�h*q��fVWVAR �<�mMx�d R e�p�bua�_DEFPROG� %�i%M�AIN TORN�O 0 RVIS�I�`�rISPL�AY�`�n�rINST_MSK  �|� �zINUSsER �tLCK)���{QUICKMEx�pO��rSCREl����+rtpsc�t)������b���_��STz�iRA�CE_CFG U=�iMt�`	nt�
?��HNL C2>�z���T{ zr @�R�d�v����������К�ITEM 2�?,� �%$1�23456789y0�%�  =<�xC�U�]�  !c�k�wp'���ns�ѯ 5����k������j� ů��鯕���A�1�C� U�o�y�󿝿I�oρ� 忥�	��-ϧ�Q��� #�5ߙ�A߽�����e� �������M���q߃� L��g��ߋ���� %�w� �[���+�Q� c���o��������3� ��{�;������ G_����/�S e.�I�m� ��=�a/ 3/������k/ /�/�/�/]/?�/�/ �/?�/u?�?�??�? 5?G?Y?�?+O�?OOaO �?mO�?�?�OO�OCO __yO+_�O�Ox_�O �_�O�_�_�_?_�_c_ u_�_o�_Wo}o�o�_ �oo)o;o�o�oqo1 C�oO�o�o�� %��[��Z���S�@��_��g  ے_� ����y
 Ï�Џ����UD1:\����q�R_GR�P 1A �� 	 @�pe�w��a���������ߟ͞� ���ّ�>�)�b�M�?�  }���y� ����ӯ������	� �Q�?�u�c���������Ϳ�	-���~o�SCB 2B{� h�e�wωϛ���Ͽ�������e�UT�ORIAL C�{��@�j�V_CONFIG D{����������O�OUT?PUT E{����������� %�7�I�[�m���� �����������%� 7�I�[�m�������� ��������!3E Wi{������ ��/ASe w������� //+/=/O/a/s/�/ �/�/�/�/��/?? '?9?K?]?o?�?�?�? �?�?�/�?�?O#O5O GOYOkO}O�O�O�O�O �O�?�O__1_C_U_ g_y_�_�_�_�_�_�O �_	oo-o?oQocouo �o�o�o�o�o�_�o );M_q�� ����yߋ���� -�?�Q�c�u������� ��Ϗ���o�)�;� M�_�q���������˟ ݟ� ��%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���
� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� �1CUgy� ������	 -?Qcu��������/�x���$/6/ !/a/ ��/�/�/�/�/�/�/ ??'?9?K?]?�? �?�?�?�?�?�?�?O #O5OGOYOkO|?�O�O �O�O�O�O�O__1_ C_U_g_xO�_�_�_�_ �_�_�_	oo-o?oQo cot_�o�o�o�o�o�o �o);M_q �o������� �%�7�I�[�m�~�� ����Ǐُ����!� 3�E�W�i�z������� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�o�~���$TX_SCR�EEN 1F8%�  �}��~���������
�� ��m&��\�n߀ߒߤ� ��-�?������"�4� F��j��ߎ����� ����_����0�B�T� f�x����������� ����>��bt ����3�W (:L^��� �����e/� 6/H/Z/l/~/�//�/��$UALRM_�MSG ?����� �/���/�/)? ?M?@?q?d?v?�?�?��?�?�?�?O�%SEoV  �-EF��"ECFG Hv����  ���@�  AuA  w Bȁ�
 O ���ŨO�O�O�O�O_�_&_8_J_\_jWQAG�RP 2I[K 0��	 �O�_� �I_BBL_NO�TE J[JT?��l�����g@�RDEFP�RO� %�+ (?%MAIN�_2m%OVoAozoeo�o�o �o�o�o�o�o@��[FKEYDAT�A 1K�ɞPp jG���_��0����z,(�����(POINT�  ]'�)�  I�RECT}@o�V�N�Dh���� CHO�ICEB���TOUCHUP׏؏� '��K�2�o���h��� ��ɟ۟���#�5���Y��y��/f�rh/gui/w�hitehome.pngd�����Ư�دꯀ{�point���0�B�T�f����  |�direc�����ƿؿ�y�/in��#�5�G�Y��k�����choic ��ϰ������������{�touchup�0�B�T�f�x���}{�arwrg� ���������߁��)� ;�M�_�q����� ���������%�7�I� [�m����������� ������3EWi {������ �/ASew� �r������/ !/(E/W/i/{/�/�/ ./�/�/�/�/??�/ /?S?e?w?�?�?�?<? �?�?�?OO+O�?OO aOsO�O�O�O8O�O�O �O__'_9_�O]_o_ �_�_�_�_F_�_�_�_ o#o5o�_Goko}o�o �o�o�oTo�o�o 1C�ogy��� �P��	��-�?� Q��u���������ϏZj�܋�u�܏��(�s��Q�c�r�,�I���A�OINT � ]���� OOK� Tß�}�NDI�RECܟ�  CHOICE�����UCHUPG�H�s� ��~�����߯�د� ��9�K�2�o�V��������ɿ��whitehom����%��7�I�X���poin��ߍϟϱ�����d�i/look}���(�:�L�^�i�indirec|Ϙߪ߼������g�choic ���� �2�D�V�h�k�touchup������������g�arwrg��"�4�F�X� j�a������������� w�0BTfx ������� ,>Pbt� �����/�(/ :/L/^/p/�//�/�/ �/�/�/ ?׿�/6?H? Z?l?~?�?�/�?�?�? �?�?O�?2ODOVOhO zO�O�O-O�O�O�O�O 
__�O@_R_d_v_�_ �_)_�_�_�_�_oo *o�_No`oro�o�o�o 7o�o�o�o&�o J\n����E ����"�4��X� j�|�������A�֏� ����0�B�яf�x� ��������O�������,�>�<L��>����u��� ��q���ͯ��,���� ��"�	�F�X�?�|�c� ������ֿ������ 0��T�f�Mϊ�qϮ� �����������,�>� ?b�t߆ߘߪ߼�˟ ������(�:�L��� p�������Y���  ��$�6�H���l�~� ����������g���  2DV��z�� ���c�
. @Rd����� ��q//*/</N/ `/��/�/�/�/�/�/ �//?&?8?J?\?n? �/�?�?�?�?�?�?{? O"O4OFOXOjO|OS� �O�O�O�O�O�OO_ 0_B_T_f_x_�__�_ �_�_�_�_o�_,o>o Poboto�oo�o�o�o �o�o�o:L^ p��#����  ���6�H�Z�l�~� ����1�Ə؏����  ���D�V�h�z����� -�ԟ���
��.� ��R�d�v�������;� Я�����*���N��`�r����������@�����@������	��+�=��,)�n�!ߒ�y϶��� �������"�	�F�-� j�|�cߠ߇����߽� ������B�T�;�x� _���O������� �,�;�P�b�t����� ����K�����( :��^p���� G�� $6H �l~����U ��/ /2/D/�h/ z/�/�/�/�/�/c/�/ 
??.?@?R?�/v?�? �?�?�?�?_?�?OO *O<ONO`O�?�O�O�O �O�O�OmO__&_8_ J_\_�O�_�_�_�_�_ �_�_��o"o4oFoXo joq_�o�o�o�o�o�o �o�o0BTfx ������� �,�>�P�b�t���� ����Ώ������(� :�L�^�p�������� ʟܟ� ����6�H� Z�l�~������Ưد ������2�D�V�h� z�����-�¿Կ��� 
�ϫ�@�R�d�vψ� ��)Ͼ��������ߴ*�`,��`���U�g�y�Q��߭߇�,���ߑ�� ��&�8��\�C��� y������������ 4�F�-�j�Q���u��� ���������_B Tfx������ ��,�Pb t���9��� //(/�L/^/p/�/ �/�/�/G/�/�/ ?? $?6?�/Z?l?~?�?�? �?C?�?�?�?O O2O DO�?hOzO�O�O�O�O QO�O�O
__._@_�O d_v_�_�_�_�_�___ �_oo*o<oNo�_ro �o�o�o�o�o[o�o &8J\3�� �����o��"� 4�F�X�j�������� ď֏�w���0�B� T�f�����������ҟ ������,�>�P�b� t��������ί�� ���(�:�L�^�p��� �����ʿܿ� Ϗ� $�6�H�Z�l�~�Ϣ� ����������ߝ�2� D�V�h�zߌ�߰��� ������
��.�@�R�d�v���qp��}�qp�����@����������,	 N�r�Y��������� ������&J\ C�g����� ��"4X?| �m�����/ �0/B/T/f/x/�/�/ +/�/�/�/�/??�/ >?P?b?t?�?�?'?�? �?�?�?OO(O�?LO ^OpO�O�O�O5O�O�O �O __$_�OH_Z_l_ ~_�_�_�_C_�_�_�_ o o2o�_Vohozo�o �o�o?o�o�o�o
 .@�odv��� �M����*�<� �`�r���������̏ �����&�8�J�Q� n���������ȟڟi� ���"�4�F�X��|� ������į֯e���� �0�B�T�f������� ����ҿ�s���,� >�P�b��ϘϪϼ� �����ρ��(�:�L� ^�p��ϔߦ߸����� ��}��$�6�H�Z�l� ~������������ �� �2�D�V�h�z�	� ������������
�������5GY1{�g,y�q�� �<#`rY� }�����/&/ /J/1/n/U/�/�/�/ �/�/�/�/ݏ"?4?F? X?j?|?���?�?�?�? �?�?O�?0OBOTOfO xO�OO�O�O�O�O�O _�O,_>_P_b_t_�_ �_'_�_�_�_�_oo �_:oLo^opo�o�o#o �o�o�o�o $�o HZl~��1� ���� ��D�V� h�z�������?�ԏ� ��
��.���R�d�v� ������;�П���� �*�<�?`�r����� ������ޯ���&� 8�J�ٯn��������� ȿW�����"�4�F� տj�|ώϠϲ����� e�����0�B�T��� xߊߜ߮�����a��� ��,�>�P�b��߆� ��������o��� (�:�L�^�������� ��������}�$6 HZl������ ��y 2DVhhzQ�|�Q�����������,�/./�/ R/9/v/�/o/�/�/�/ �/�/?�/*?<?#?`? G?�?�?}?�?�?�?�? OO�?8OO\OnOM� �O�O�O�O�O�O�_ "_4_F_X_j_|__�_ �_�_�_�_�_�_o0o BoTofoxoo�o�o�o �o�o�o�o,>P bt����� ���(�:�L�^�p� ����#���ʏ܏� � ���6�H�Z�l�~��� ���Ɵ؟���� � ��D�V�h�z�����-� ¯ԯ���
����@� R�d�v��������Oп �����*�1�N�`� rτϖϨϺ�I����� ��&�8���\�n߀� �ߤ߶�E�������� "�4�F���j�|��� ����S�������0� B���f�x��������� ��a���,>P ��t�����] �(:L^� ������k / /$/6/H/Z/�~/�/@�/�/�/�/�/���+��������?'?9=?[?m?G6, YO�?QO�?�?�?�?�? OO@ORO9OvO]O�O �O�O�O�O�O_�O*_ _N_5_r_�_k_�_�_ �_�_��oo&o8oJo \ok/�o�o�o�o�o�o �o{o"4FXj �o������w ��0�B�T�f�x�� ������ҏ������ ,�>�P�b�t������ ��Ο������(�:� L�^�p��������ʯ ܯ� ���$�6�H�Z� l�~������ƿؿ� ��ϝ�2�D�V�h�z� ��ϰ���������
� ��_@�R�d�v߈ߚ� �Ͼ���������*� ��N�`�r����7� ��������&���J� \�n���������E��� ����"4��Xj |���A��� 0B�fx� ���O��// ,/>/�b/t/�/�/�/ �/�/]/�/??(?:? L?�/p?�?�?�?�?�? Y?�? OO$O6OHOZO��$UI_INU�SER  ����{A��  [O_O_M�ENHIST 1�L{E  �(�@3�(/�SOFTPART�/GENLINK�?current�=menupage,153,1�O0__1_C_�'�O�N�71�@BARRA�_ESTEIRA �O�_�_�_�3)X_�E�edit�BMAI=N�QACE0�_o�.o@o�90�_�^PE�GA_TORNO,13Lo�o�o�o�8s� ao�M962o�-?Q�o�oq36
����dv�A48,2�%�7� I�[����O����Ǐُ�3���0�A��� �"�4�F�X�j�m��� ������ȟڟ�{�� "�4�F�X�j������� ��į֯�w���0� B�T�f�x�������� ҿ������,�>�P� b�t�ϘϪϼ����� ����(�:�L�^�p� �߅�#߸������� � ��6�H�Z�l�~�� ������������� ��D�V�h�z�����-� ��������
��@ Rdv��);� ��*�N` r������� //&/8/�\/n/�/ �/�/�/E/�/�/�/? "?4?F?�/j?|?�?�? �?�?S?�?�?OO0O BO�?fOxO�O�O�O�O �OaO�O__,_>_P_ ;t_�_�_�_�_�_�_ �Ooo(o:oLo^o�_ �o�o�o�o�o�oko  $6HZl�o� �����y� � 2�D�V�h�������� ԏ������.�@��R�d�v�aX�$UI�_PANEDAT�A 1N������  	��}  frh�/gui��dev�0.stm ?_�width=0&�_height=�10ԐÐice=�TP&_line�s=15&_columns=4Ԑ�font=24&�_page=wh�oleÐ��\V) � rim#�L�   ��c�u���������$� ϯ�گ���;�M�4� q�X�������˿������%�\V� ��   
 � ���]���cgtp/flexÐ(Ǒ̟ޛ2�3t����1
�doubÐ2/�-�ual����_� �"�4�F�X�j�ώ� u߲��߫������� �B�)�f�M�������3�E�  �������*�<� N�`�����Ϩ����� ����i�&8\ C��y���� ��4Xj=���������� � /S$/��H/Z/l/ ~/�/�/	/�/�/�/�/ �/ ?2??V?=?z?a? �?�?�?�?�?�?
O} �@OROdOvO�O�O�? �O1/�O�O__*_<_ N_�Or_Y_�_}_�_�_ �_�_�_o&ooJo1o no�ogo�oO)O�o�o �o"4�oXj�O ������O� �0�B�)�f�M����� ���������ݏ�� >��o�o��������� Ο��3��w(�:�L� ^�p���韦�����ܯ ï ����6��Z�A� ~���w�����ؿ�]� o� �2�D�V�h�z�Ϳ �����������
�� .ߕ�R�9�v�]ߚ߬� ���߷������*��@N�`�G����	����@���������"�)�� G���6�s��������� ��4�������K 2oV���������#������$UI_POST�YPE  ��� 	 �/�UQUICK�MEN  d�s�WRESTO�RE 1O��  ���� /#���m +/T/f/x/�/�/?/�/ �/�/�/?�/,?>?P? b?t?/�?�?�??�? �?OO(O�?LO^OpO �O�O�OIO�O�O�O _ _�?_1_C_�O~_�_ �_�_�_i_�_�_o o 2o�_Vohozo�o�oI_ So�o�oAo�o.@ Rd����� s���*�<��oI� [�m������̏ޏ�� ���&�8�J�\�n���������ȟڟ�SC�RE�?��u1sc�uU2�3�4�5��6�7�8��T;AT`� ��MUSER�����Sks���3��4��U5��6��7��8���UNDO_CFG� Pd����UP�DX�����None���_I�NFO 1Q�<��0%��W��� E���i��������� տ���:�L�/�pς��eϦύ)�OFFS�ET Td@� ��{������	��-� Z�Q�cߐ߇ߙ��ϝ� ������ ��)�V�M�_�q�۹�����
����t��)�WOR/K U4������A�S��ψ�UFRAME  ���&��RTOL_ABRqT��$���ENB��~��GRP 1V���Cz  A� ��+=Oa s�����U����~��MSK  ��<���N��%4���%��)��_EVN������>�2W���
 h��U�EV��!td:�\event_u�ser\-�C7ȍ��}�F��SP���spotw�eld�!C6 ����!� Z/�/:'�H/~/l/�/ �/�/�/-?�/Q?�/?  ?�?D?�?h?z?�?O �?)O�?�?OqO`O�O @ORO�OvO�O_�O�O@7_�O[__Z]W+�32X����8V_�_�_ �_�_o�_,o>o obotoOo�o�o�o�o �o�o�o:L'�p�]����$�VARS_CON�FI�Y�� FP�{���|CCRG��\��>�{��t�D� BH� p,k�a�C�� ��}��?���C,&Q=��mͩ�A �MR;2b���	}��	��@�%1: �SC130EF2� *����{�����,X� �5}������A@k�C�F� 	w�Q�[���|��� �������T�����\�ϟ �\� B���;�e�@�ǟ `�����S�����̯�� �ۯ�&�}��\�G��Y���E���ȿ�TCC�c
�������M�pGF�pgd���-�2345?6789017�?��ׁ$���4�v�N m�� ��϶�BW������i�}�:�o=LA�څ�6�@�6�Ϳ�Z���i�7����(�� W���-�]�X�jĈߚ� �ϳϹ��������� %�7�I�r�m�ߨ�� �����������8�3� E�W������}����� ��������/�A�S�xe�w��MODE���t �RSLTg e�|k�%"z� ���;�1��d���`��SELEC���c��	IA_[WO�Pf ��� W,		�������G�P ������RTSYONCSE� ��$��	#WINURL 3?*ـ�;\/�n/�/�/�/�/�uISIONTMOU����A# ��%�g�Sۣ�SۥP��� FR:\~�#\DATA\�/� �� MC�6LOG?   oUD16EX@?�\�' B@ ����2T1  a�briel_Fariak?P5�?�?������ n6 � ���GV�2\�� -��5�� C  ��Z�@U058TRAINj?��*B�{Rd_Cp��D #`{2��'$�":��h#� (�kI �Mw��O�O�O�O�O1_ _U_C_]_g_y_�_�_\�_�(STA� i�@�@�o o2oI8$>o\bo�%_GE�j#�;�~@ �
�\�|�btgHOMIN�_kSۮ��`�2(,,��CWǖBve�JMPERR 2=l#�
  ��I: ��"�4Fwj| ��������l�&%S_g0RE鰹m�^۴LEXdn��1-ehoVM�PHASE  �e׃BޱOFF� _ENB  ޢ$VP2�$oS�ۯ��x�c C�;�@ �a;���?Gs33'D*AA���]� ��0ޱ�`r�}�XC��܅���� ��[�6�������6��]���>VYD-۟�E B�[��t\16���+FV���W��5d����� ,�>�'Es���W�I�ǟ��� ��I���� �9�k�ɯ;������� ׯɿ3�տ����C�8� g�Yϋ��ϯ���ϱ� ������-�"�Q�c�u� jߙ�?��ϗߩ߻��� �u���M�B�T��u� �߁��������� 7�,�[�m��]�k�}� ���������!�E� ����CUg���! ���� /!�- WQ������ c	//)/?/M'�s�TD_FILTuE�`s�k �x2�`����/�/�/�/ �/	??-???Q?�6�/ ~?�?�?�?�?�?�?�?�O OoiSHIFTMENU 1t}<5�%5�~O)�\O �O�O�O�O�O�O�O'_ �O_6_o_F_X_�_|_��_�_�_	LIV�E/SNAP�S?vsfliv���_��z`ION �ҀU
`bmenu &o+o�_�o�oV"<E�uz��4IMO�v����zq�WAIT�DINEND  a�ec��b�fOKوNOUT�hSD�yTIMdu��o|G�}#�{C�z�b�z�xRELE���ڋxTM�{�d=��c_ACT`و���x_DATA �wz���%  E�GA_BARRA�_ESTEIRAx�o6Ex�RDIS
`~E��$XVR�a�x�n�$ZAB�C_GRP 1yvz��� ,��2̏.MZD��CSKCH�`z���aP@��h@�IP�b{'���şן�[��MPCF_G 1|'���0�r�8�d�� �}'�(�p�s�� 	(���  �<l0  ���?�A�M\����5���������|2MP�����A  %Cj�_�D���1w��?Ý���{b�?7N��b���=.I ������ɯۯ������o���w���� �/��3���7?�lB� ˿ݸ ĸ+��	��1�?�i���'�9�0?�Q���	��`~����_CY�LIND~!�� Р ,(  *.�?ݧ+�h�O���s� �������� (�	�x�-��&�c�� ��������j�P�� ��)��~�_�q��� �s2�'��� �&� ���������&���I��cA���S�PHERE 2��������� �A�T/A��e ������/ N`=/�a/H/Z/�/`��/�/�/��ZZ� ��f