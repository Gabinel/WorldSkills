��   T�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ������DMR_SHF�ERR_T  � $OFF�SET   w	  /GRP:�� $MA���R_DONE � $OT_M�INUSJ  	�sPLzdCOU=NJ$REFj��PO{��I$�BCKLSH_S�IG�EACH�MSTj�SPC��
�MOVn ~A�DAPT_INE�RJ FRIC�COL_P,MGRAV�� �HISIDSP|k�HIFT_7 -O �Nm��MCH� S�AR�M_PARAO� dcANGo zy2�CLDE7��CALIBD~n$GEAR�=2� RING���<$]_d�REyL3� 1 N ��CLo: �� �AX{  o$PS_�TI����TIME z�J� _CMD���"FB�VA �&C�L_OV�� FR�MZ�$DEDXv�$NA� %�OCURL�W����TCK�%�F�MSV�M_LIF	��'8�3:c$�-9_09:_ ��=�%3d6W� �">�PCCOM���FB� M�0�MAL_�ECI��P:!o"DTYkR�_|"�5:#�1END��4��o1 el5M�P PL� �W ��STA>:#TRQ_M���� KNiFS� uHY�sJ� hGI�JI�JI�D �$�ASS�> ����A������@VERSI�� �G  �0��AIRTU�AL�O�AS 1~�H ���N ��\_G_�_k_ �_�_�_�_�_�_�_���Po�DBo0l�YH�v ��� ��"��
 9d���A/o�o+oUl�o@�o�o�o�o�k;�Ar*gyd���d�������=L̙���?����@�=�b�t����������Ώ�����(�{ �US�a�K����D  2���ğ֟���@��0�B�T���<�� ~�������Ưد����� �2�D���Pr�( �x����������� Ͽ���>�)�b�Mϰ��qϖϼ��$4 �12\���M{�ֽJ���K��БU�2[V,��lP��d��E��f�HZR"E���~;d�;<�>;���A���Aߚ�h�z�e� ��9�K߅���߈��� �9�$�]�o��X�L�X�fqX����� ���T���@P������'���%���345678901G�O�t�x�q���m� ����������D� }���z�H��lZ| �����.�� 2 Vh���� n@���/r� U/���//�/�/�/ �/8/	??n/�/N?<? r?`?�?�?�/�?"?4? �?�?O8O&O\O�?�? �O�?�?�OFO�O�O�O "_xOI_[_�O_�_|_ �_�_�_�_>_ob_t_ �_�_Boxofo�o�_o �o(o:o�o,< b�o���oP�� ���(�~O��� .� �������܏2�D� �h�z�H�Əl�Z�|� ����ɟ۟.������ 2� �V�h�������� n�@�¯����r��� U�������������� �8�	��n�пN�<� r�`ϖϨ�����"�4� �π��8�&�\�n�}�p�ϕ����60�����9��$PLCL�_GRP 1S��� D�?�  ��� ;��_�J��n��� ���������%��