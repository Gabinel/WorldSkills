��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@  &��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	�>&USRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  w0�aIRTs1�	o`'2 L1��L1��R�	 �,��?���a�1`�b�ba ����� _�  ?����
 ��a�o�o 1CU �oz �����c�
� �.�@�R��v����� ����Џ�q���*� <�N�`�������� ̟ޟm���&�8�J� \�n���������ȯگ �{��"�4�F�X�j� ��������Ŀֿ����`TPTX������/�` �sȄ�$/so�ftpart/g�enlink?h�elp=/md/�tpmenu.dg���ϨϺ��υ��� ��&�8�J���n߀� �ߤ߶���W������ "�4�F�X���|��ﰲ��������ar�f�b�� ($p�-����T�?�x��� a�a��c���c����l��c�g���a�a�a��ah��a2�h�	.f���������8�a���`  ���f >ep��h%#h�F�bc Xc�B� 1)hR �\ _�� �REG VED�]���whol�emod.htm��	singl	�doub t�rip8browsQ���� �u���//@/����dev.Esl�/3� 1�,	t�/_�/;/i/? ?/?�/S?e?w?�?�?�?� ��?�?O O%O7OIO[OmOO�E 2P�?�O�O�O�O�O_ �E�	�?�?;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omooM' �o�o�o�o�o�o +=Oas��� ������?>�P� b�t���������Ώ�� �O�����L�^�_ '_�������ş�� ���6�1�C�U�~�y� ����Ư��ӯ�o�� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�-��ϬϾ��� ������*�<�7�`� r�A�Sߨߺ�q���i� ����!�J�E�W�i� ������������� "��/���O�I�w��� ������������ +=Oas��� ����,>P bt���߼�� �//�����^/Y/ k/}/�/�/�/�/�/�/ �/?6?1?C?U?~?y? �?Y��?�?�?�?�?	O O-O?OQOcOuO�O�O �O�O�O�O�O__� R_d_v_�_�_�_�_�_ �_�_�o*o�_o`o�ro�j�$UI_T�OPMENU 1�K`�aR� 
d�a*Q)�*defaul�t5_]*le�vel0 * [	G �o�0�o�'rtpio[2�3]�8tpst[1[x)w9�o	��=h58E01?_l.png��6?menu5�y�p��13�z��z	�4���q��]����� ����̏ޏ)Rr����+�=�O�a���pr�im=�page,1422,1h� ����şן�����1�C�U�g���|�c?lass,5p������ɯۯ�����13��*�<�N�`�r���|�53������ҿ(�����|�8��1� C�U�g�y����ϯ���������"Y�`�a�o /��m!ηq�Y��av�tyl}Tfqmf[�0nl�	��c[1364[w��59[x�q�G�y��tC8�|�2 9��o�%�1���{�� m��!�����0�B� ��f�x���������o���80��'9K~���2P��� ��\��'9 K������������1��/$/6/�H/Z/U�|�ainedi'ߑ/�/�/�/��/P�confi�g=single}&|�wintp�� �/$?6?H?Z?	�ߐ?|?ٷ�gl[57��@�q��?�;gp�08�݂�07I�?F��F2JO[6�:�?)O�O�xl �� �4s�x �O���$��`�o�H_ Z_l_~_�_�_Q��_�_ �_�_o o�_DoVoho�zo�o�o�o�!;�$d�oub5o��13���&dual�i38��,4�o&�o9�o�n�o�a8�� �Ao����&�8�
�%3L=}!��o�b8@���������z� ��(�:��+:T��i48,2o��b{����ʟ {?�;�M� sc���;���s�� �}���e�u��X��@�F7L���`�O��2�4h�z�6e�u7���� �ｿϿ���̏�27��G�Y�k�}Ϗ� �0�s��������
�!�1�M�_�q� �ߕ����������� ��7�I�[�m��� ������������!�����6(�]�o��������$��746�����)�C�ߟT��	TPTX[209�<Aw2IHJ���Bw1H�]H���(��02��A0#��[Ttv`��O�L#_�0� \��5S�[�treevie�w3v�3��~�381,26M/_/q/ 0�/�/�/�/�/�/~/ ?%?7?I?[?m?�o/�(��o5%���?�?�?��A�?\1~��?8"2 ��eOwO�?�?(}�LE K��O�O_�O��8@�O NOa_s_�_��6_d� E_�_�_�_oV�#_�� �_�Sooo�o�oB�o �o��oA�oq +=Oas��o� ������(�9� ��Q�x���������ҏ ?����,�>�P�ߏ t���������Ο]��� ��(�:�L�^�ퟂ� ������ʯܯk� �� $�6�H�Z��l����� ��ƿؿ�y�� �2� D�V�h����Ϟϰ��� ���ϕo�o��o@ߧ E�c�u߇ߙ߽߬��� ��O����)�<�M�_� q���W�������� �&�8���\�n����� ����E�������" 4��Xj|��� �S��0B �fx����O ��//,/>/P/� t/�/�/�/�/�/]/�/ ??(?:?L?��߂? 1ߦ?���?�?�?�? O$O5OGO�?SO}O�O �O�O�O�O�O�O��2_ D_V_h_z_�_�_�/�_ �_�_�_
oo�_@oRo dovo�o�o)o�o�o�o �o*�oN`r ���7���� �&��J�\�n����� ����E�ڏ����"� 4�ÏX�j�|������� a?s?蟗?�sO_/� A�S�e�w�������� �������,�=�O� a�#_������ο�� =��(�:�L�^�pς� Ϧϸ������� ߏ� $�6�H�Z�l�~�ߐ� ������������2� D�V�h�z������ ������
����@�R� d�v�����)����������ƚԔ*d?efault%���*level8��ٯw���? �tpst[1]��	�y�tpi�o[23���u����J\me�nu7_l.pn5g_|13���5�{�y4�u6���//'/9/K/ ]/���/�/�/�/�/�/ j/�/?#?5?G?Y?k?~�"prim=|�page,74,1p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_0f_x_{?�218�?�_@�_�_�_�__B6o�9oKo]ooo�o`�$�UI_USERV?IEW 1֑֑�R 
���o��o�o[m�o'9K]  �����l�� �#�5��oB�T�f�� ����ŏ׏鏌��� 1�C�U�g�
������� ��ӟ~�����v�?� Q�c�u���*�����ϯ �󯖯�)�;�M�_� 
��~������ݿ� ��%�ȿI�[�m�� ��4ϵ��������Ϩ� 
��.ߠ�i�{ߍߟ� ��T���������/� ��S�e�w���Fߨ� ����>���+�=�O� ��s���������^��� ��'����FX ��|������ #5GY�}� ���p���h 1/C/U/g/y//�/�/ �/�/�/�/�/?-??? Q?c?/p?�?�??�? �?�?OO�?;OMO_O qO�O&O�O�O�O�O�O �?�O_ _�OD_m__ �_�_�_X_�_�_�_o !o�_EoWoio{o�o0h