��   g�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����BIN_CFG_�TX 	$EN�TRIES  �$Q0FP?N�G1F1O2F2�OPz ?CNET�G���DHCP�_CTRL. � 0 7 ABL�E? $IPUS~�RETRAT��$SETHOS�T��NSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM�� !� FT�� @� LOG_�8	,CMO>$�DNLD_FIL�TER�SUBDIRCAPC��\8 . 4� H�{ADDRTYPz�H NGTH�̉��z +LS�q D $R�OBOTIG �P�EER�� MAS�K�MRU~OM�GDEV��PI�NFO�  {$$$TI ��RCM+T A$( </�QSIZ�!�S� TATUS_�%$MAILSE�RV $PLA�N� <$LIN><$CLU���<$TO�P$C�C�&FR�&YJE�C|!Z%ENB �� ALAR:!BF�TP,�#,V8 }S��$VAR�)�M�ON�&���&A7PPL�&PA� �%���'POR�Y#_|�!�"ALERT�&�i2URL }>Z3ATTAC��0�ERR_THRO�U3US�9H!�8� CqH- c%�4MAX?wWS_|1��1'MOD��1I�  ��1o (�1PWD  � LA��0��ND�1TRYFD�ELA-C�0G'AE�RSI��1Q'RO.BICLK_HM 0Q'ί XML+ 3SG�FRMU3T� !O�UU3 G_�-COAP1�F33�AQ'C[2�%�B_AU�� 9 �R�!UPDb&P�COU{!�CFO 2 
$V*W8�@c%ACC_HYQ�SNA�UMMY�1oW2"$DM*�  $DIS��SM	 !l5�o!�"%Q7�IDZP�%� �VR�0z�UP� _DLVS'PAR��QN,#�
3 �_�R!_W�I�CTZ_IND9E�3^`OFF� ~URmiD�)c�   t Z!N`MON��cD�.�bHOUU#E%A�f��a�f�a�fLOCAܗ #$NS0H_[HE���@I��/  d8`ARP�H&�_IPF�W�_* O�F``QF�AsD90�VHO_�� 5R42PSWq?�wTEL� P����90WORjAXQE� LVt�[R2�ICE���p� �$cs  O����q��
���
�p�PS�A�w[# 0�	�Iz0�AL��' �
���F����!�p��i��$� 2Q��P���������� Q���!�q�����$� _FLTR � �\� ��
��������$Q��2��7rSH`D +1Q� P㏙�f���ş��韬�� П1���=��f���N� ��r�ӯ�������ޯ �Q��u�8���\��� ����󿶿�ڿ;��� _�"�XϕτϹ�|��� ��������6�[�� �Bߣ�f��ߊ��߮� ��!���E��i�,�� P�b���������� /���(�e�T���L���l��z _LUA1�_x!1.��0���p���1��p�25c5.0��r��n���2����d %7I[3e��� ����[4���T'9[5U��� {���[6���@D �//)/s��Q�ȁMA��M?A� ����� Q� ��u.<�/?&?�/J?\? n?A?�?�?m�P�?�? �?�?�?O.O@OROOvO�O�Ou.kOl�q���O�L
ZDT ?StatusZO�O�5_G_Y_n�}iR�Connect:� irc{T//alert^�_�_�_ �_mW#_oo,o>oPo�bot�^�d~2g���go�o�o�o�o�o�o 	-?Qcul��$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5_3e036�`(�_��_���"�p�1!W��(��"S��J�E�� X��tQ���,$���W���ˏ�� �֏��%��I�0�m� �f�����ǟ��������!��u�R������ DM_�!�����SMTP_C?TRL 	����%����DF���ۯ�t�ʯ��'��Lz�N���!
j��y�q�>u����Ԙ��#�L�USTOM �j������  |���$TCPIPd��j��H�%�"�E�L�����!���H�!TP��j�?rj3_tp�b;����i�!KCL�G�L�i���5�!C�RT�ϔ����"u�?!CONS��M��[�ib_smo	n����