��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@)8&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	�>&USRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  w0�aIRTs1�	o`'2 L1��L1��R�	 %,��?���a1`#�b�d~a���c��� � � �o��
 ��a�o�o1CU �oz���� �c�
��.�@�R� �v���������Џ� q���*�<�N�`�� ��������̟ޟm�� �&�8�J�\�n����� ����ȯگ�{��"� 4�F�X�j����������Ŀֿ���`/TPTX������/�` sȄ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ� ���υ�����&�8� J���n߀ߒߤ߶��� W������"�4�F�X� ��|�����������a�`��b�� ($p�-����T�?�x���a�a��cH���g��l��k
����a��h�ah��a2�h�	f����������`���`�  ���f ep���h#h�F�bc Xc�B 1~)hR \ �_�b REG VED]����wholemo�d.htm�	si�ngl	dou�b trip�8brows Q�����u� ��//@/����dev.slh�/3� 1�,	t�/ _�/;/i/??/?�/�S?e?w?�?�?�?� ��?�?OO%O7O`IO[OmOO�E @�? �O�O�O�O�O_�F�	 �?�?;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omooM'�o�o �o�o�o�o+= Oas����� ����?>�P�b�t� ��������Ώ���O� ����L�^�_'_� ������ş����� 6�1�C�U�~�y����� Ư��ӯ�o���-� ?�Q�c�u��������� Ͽ����)�;�M� _�-��ϬϾ������� ��*�<�7�`�r�A� Sߨߺ�q���i���� �!�J�E�W�i��� �����������"�� /���O�I�w������� ��������+= Oas������ �,>Pbt ���߼���/ /�����^/Y/k/}/ �/�/�/�/�/�/�/? 6?1?C?U?~?y?�?Y� �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__�R_d_ v_�_�_�_�_�_�_�_ �o*o�_o`oro�j��$UI_TOP�MENU 1�K`�aR �
d�a*Q)*default5_�]*leve�l0 * [	 �o�0�o'r�tpio[23]��8tpst[1�[x)w9�o	�=�h58E01_l�.png��6m�enu5�y�p�1!3�z��z	�4���q��]��������� ̏ޏ)Rr���+�=��O�a���prim�=�page,1422,1h����� şן����1�C��U�g���|�class,5p�����ɯhۯ�����13��@*�<�N�`�r���|�53������ҿ���
��|�8��1�C�U� g�y����ϯ���������"Y�`�a�o/��m�!ηq�Y��avtyxl}Tfqmf[0n�l�	��c[164[w��59[x�qG�y�&�tC8�|�29�� o�%�1���{��m�� !�����0�B���f��x���������o���80��'9K~���2P����� \��'9K� �����������1��/$/6/H/Z/�U�|�ainedi'ߑ/�/�/�/�/P��config=single&|�wintp���/$? 6?H?Z?	�ߐ??ٷ�gl[57�ٳqߐ�?�;gp�08�ݲ07�I�?F��F2JO[6�:�?)O�O�x �� �4s�x�O�� �$��`�o�H_Z_l_ ~_�_�_Q��_�_�_�_ o o�_DoVohozo�o�o�o�!;�$dou�b5o��13��&odual�i38��C,4�o&�o9�o �n�o�a8���Ao�����&�8��%3BL=}!��o�b8@� ��������z����(�:��+:T��i48,2o��b{����ʟ {?�;�M�sc���;���s�� �}����e�u��X��@�F7 L���`�O��2�h�z�6e�u7�����ｿ�Ͽ���̏�27 ��G�Y�k�}Ϗ��0Ās���������!�1�M�_�q߃ߕ� ������������ 7�I�[�m����� ���������!�����6(�]�o��������$��746������)�C�ߟT�	TPTX[209�<Aw2IHJ���Bw1H�]H����
�02��A#��[Ttv`��O�L#_��0� \��5S[�treeview3�v�3��~�381,26M/_/q/0�/ �/�/�/�/�/~/?%? 7?I?[?m?�o/(��o`5%���?�?�?�A�?"\1~��?8"2��eO wO�?�?(}�LEK��O �O_�O��8@�ONOa_s_�_��6_d�E_�_ �_�_oV�#_���_�S ooo�o�oB�o�o� �oA�oq+= Oas��o��� ����(�9���Q� x���������ҏ?�� ��,�>�P�ߏt��� ������Ο]����� (�:�L�^�ퟂ����� ��ʯܯk� ��$�6� H�Z��l�������ƿ ؿ�y�� �2�D�V� h����Ϟϰ������� �o�o��o@ߧE�c� u߇ߙ߽߬�����O� ���)�<�M�_�q�� ��W���������&� 8���\�n��������� E�������"4�� Xj|����S ��0B�f x����O�� //,/>/P/�t/�/ �/�/�/�/]/�/?? (?:?L?��߂?1ߦ? ���?�?�?�?O$O 5OGO�?SO}O�O�O�O �O�O�O�O��2_D_V_ h_z_�_�_�/�_�_�_ �_
oo�_@oRodovo �o�o)o�o�o�o�o *�oN`r�� �7�����&� �J�\�n��������� E�ڏ����"�4�Ï X�j�|�������a?s? 蟗?�sO_/�A�S� e�w����������� ����,�=�O�a�#_ ������ο��=�� (�:�L�^�pς�Ϧ� �������� ߏ�$�6� H�Z�l�~�ߐߴ��� ��������2�D�V� h�z���������� ��
����@�R�d�v� ����)����������ƚԔ*def�ault%��*?level8�ٯ�w���? t?pst[1]�	��y�tpio[#23���u����J\menu7_l.png_M|13��5�h{�y4�u6� ��//'/9/K/]/�� �/�/�/�/�/�/j/�/�?#?5?G?Y?k?�"�prim=|page,74,1p?@�?�?�?�?�?�"�6�class,13 �?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo�]ooo�o`�$UI�_USERVIE�W 1֑֑�R 
�A��o��o�o[m�o '9K] �� ���l���#� 5��oB�T�f������ ŏ׏鏌���1�C� U�g�
���������ӟ ~�����v�?�Q�c� u���*�����ϯ�� ���)�;�M�_�
�� ~������ݿ��� %�ȿI�[�m�ϑ�4� ���������Ϩ�
�� .ߠ�i�{ߍߟ߱�T� ��������/���S� e�w���Fߨ���� >���+�=�O���s� ��������^����� '����FX��| ������# 5GY�}��� �p���h1/C/ U/g/y//�/�/�/�/ �/�/�/?-???Q?c? /p?�?�??�?�?�? OO�?;OMO_OqO�O &O�O�O�O�O�O�?�O _ _�OD_m__�_�_ �_X_�_�_�_o!o�_ EoWoio{o�o0h