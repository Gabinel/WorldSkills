��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ��!PCOUPLE�,   $�!PPV1CES C G�1�!�� A> �1	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q�RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Nb_OPT�2 �� ELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1� UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t���MO� �sE 	� [M�s��2�wREV�BILF��1XI� %�R 7 � OD}`j��$NO`M��!b�x�/��"u�� ����4AX��@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC���a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���OR BIGALwLOW� (KtD2�2�@VAR5�d!�A}#BL[@S �� ,KJqM�H`S�pZ@M_O]z����CFd XF�0GR@��M��NFLI���;@U�IRE�84�"� SgWIT=$/0_No`�S�"CFd0M�� �#PEED���!�%`���p3`J3tV�&$E�..p�`L��ELBOF � �m��m�p/0��CP�� F�B�����1��r@1J1E_y_T>!Բ�`���g���G� �>0WARNMxp�dp�%`�V`NST� �COR-rFL{TR�TRAT �T�`� $ACC�qM�� R�r$OcRI�.&ӧRT�sSFg�0CHGV0I�p�T��PA�I{�T�!��� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8��9/C���x@�2w @� TRQ���$%f��ր����_�U������Oc <� ����Ȩ3�2^��LLECM�-�MULTIV4�"$���A
2q�CHILDh>�
1��Oz@T_1b�  4� STAY2�b4�=@�)2�4����@�� | 9$��T�A�I`�LE��eTO���E��EXT���ᗑ�B�᎞22�0>���@��1b.'��B 9�A�K�  �"K� /%�a��R���?s��?�O�!M��;A�֗�M8�� 	�  =�I�" L�0[�� �R�pA��$JOB`B���������IGI�# dӀ����R� -'r��A�ҧ_��`�n�b$ tӀFL6��BNG�A��TBA � ϑ�!��
/1�À �0���R0�P/p ,����%�|���Bq@W�
2JW�_RH�CZJZ�_zJ?�D/5C�	�ӧ���@��;�Rd&A������ȯ�qGӨ�g@NHANC��$LG/��a2qӐ� ـ�@��A�p� ���aR���>$x��?#DB��?#RA�c?#AZ�t@�(.�����`FCT����_F࠳`�SM��!I�+lA�% ` �` ���$/�/�@���[�a��M�0�\��`��أHK��A�Es@͐�!�"W��Nz� SbXYZW�`$�"����6	�������'  . I�I��2�(p�STD�_C�t�1QA��U+STڒU�)#�0U�[�%?IO1���� _Up�q�* 1\��=�#AORzs8B�p;�]��`O6  RSY�G�0�q^EUp� H`G�� ��]�@P_XWORK�+^�?$SKP_�p��DB�TR�p , �=�`����Z �m�OD3��a _C`"�;b�C� �GPL:c�a�tőS�D�W�3Bb����P�.��  @�!�-�B APR��
�qDJa3��. /��u�������LuY/$�_����0�_��/ �PC�1�_����~�EG�]� �2�_��I�
!.��R3�H $C��7.$L8c/$uSނ�z IkINE�WA_D1%�ROyp���ŀ����q�c7 t@�fP�A���RETUR�N�b��MMR"U���I�CRg`EWM�@�SIGNZ�A� ���e� 0{$P'�1$P� &m�2p�p'tm�+pD�@ �'�bdNa|)r�GO_AW ���@ؑB1@CYSd�(�CYI�4��B�`1w�qu��t2�z2�vN�}��E}s�DEVIs` 5� P $��RB���I�wPk��IG_BY���"�T7Q��tHNDG�Q6� H4��1�w��$DSBLC��o��v�g@��TPqL��70O�f@]���FB���FEra8�ׂ�t}s��
�8> i�T1?���MCS���fD �ւ
[2H� W��EE����%F��Ů@q����9� T�p��x�NK_QN:�����U��L�wKHA�vZ��~�2����P~r�q7: �N=MDLn���9�� ��ٱh����!e����J��~�+���� ,�N�D����3��Ւ8G!aqSLAd�7w;  ��INP���"�����}q_ �4<j�06`C� NU��W  D�Lק��SSH!�7=M��q���ܢӢ��������>P +$ٰ�٢��^��^�,�Y�FI B\��� ���'A	'AWl�'NTV��]�V~�X�SKI�#T���a�Hۺ�T1J�3:3_�P��SAFN���_�SV�EXCLUT��N@�DV@L���@�Y����S�HI_yV
0\2PPLYP�Ro�HIM�T�n�_�MLX��pVRF�Y_�Cl�M��IOC�UC_� ���2�O�q�LS�0v�JFT4Q�����J�@P�E$�t��A��CNFt�6եu��pm�4ACHD�o���l���AFC CPl�V�TQsP?�� �� 3?`�@TA�@�0.L@ ��N��]�' @����T��T!� S���h�e@{RA� DO�� w2L���!n��_1�B#�H!�̔�΀K���B�2��MARGIr�$����A ���_SGNE�C;
$�`�a^aR0��3���  B��B��ANNUN�P?���uCN@�`%0����� X���BEFc@I�RD @Q�F���4OT�`�sFT�HR,Qh��CQ0�M��NI|R!E�����AW����DAY=CLOAD��t;T|�<S5}�EF_F_AXI��F`�1QO3O��S�@_�RTRQE�G�����0RQj�Evp ���F�0f�R�0 �t MP�E><� H 0�``œ^�`Ds�DU�`����BCAr� �I?�`N ErID?LE_PWRI\4V!n0V�wV_[ ꐾ� �DIAG�5J�� 1$V�`SE�3TQl�e��0Pl�^E_��j��VE� �0SW�H�q(� C2�G�n�OHxPPLHk�IRAl�B�@ �[��a�bk��w3��O � ��v��I��0 �pRQDWf�MS-�%AX{<6j�LIFE�@�&�MQy�NH!Q%��$F#C����CB0��mpN$�Y @D1FL�Al���OV0]&H�E��l�SUPPO$�@u�y��@_�$�冀!_X83�$gq�'Z�*W�*B1�'T�#`�fk2XZáj�Y2D8ECY`T@�`N����f� �C�k�̒�ICTA�K `�pCACH�ӫ�3з���I��bNӰUFFI� \��@���;T��<S6CQ�����DMSW�5L �8	�KEYIMAG�cTMLa��*Ax��&E���a�rOCVI�ER-aM ��B�GL����y�?� Q	��П4N�:�ST�!�BP�D�,P�D��D��@EM�AI䐔a��sPs�FAUL|RObB�c��� spUʰ�`X DT�'`E�P< $dS�S[ � ITw��BUF�7y��7�tN�[�LSUB1T�C�x�o�R�tRSAV |U>R'c2�\�WT����P�T�*`Sn�_01PbU���YOT�bK�
�P��M��d���W#AX��2��X1P�ְS_GH#
�pYN�_���Q <��D���0���M�*� T�F�`|�\�{DI��EDT_P$ɰ:�R��b�GRQM�&��Jq�a�1׀��F�s� S (�S�VqpB��4�_�fa�u�b��T� ��@���B�SC_R]1IKU'r��$t���R"A#u�H�aDSPd:FrP�lyIM|S as�qz��a� U>w� 4<1%sM�@IP��s��0`tTHb0ЃTr2��T`asHS�cCsGBSCʴq0� V������S�_D��CONVE�G���b0$^v1PFHy�dCs�`�&aVSC���sM�ERg��aFBCM�Pg��`ET[� mUBFU� DU%Pb�D�:12�CDWy�p�P�C��R��6�:�AV� ��� ���P�ъ�C�����w������`��WH *�LƠ�Cc�W��� �Y�賂��р�q�@|���A��7}��8}�9}�H ���1���1��1��1��1�ʚ1ך1�1�2R��2����2��2��U2��2ʚ2ך2�U2�3��3��3�����3��3��3ʚ3*ך3�3�4���A'EXT[�X[b�H ``t&``z�k`˷$�����FDR�YTPV��RK"	��.K"REM*F��]"�OVM:s/�A8�T7ROV8�DT�PX�MXg�IN8ɉ W�N�INDv�["
���`K ^`G1a�a��@�Q%7Da�RIVx��u"]"GEAR:qKIO.K(�[$N�`����,(�F@� \#Z�_MCM<0K! ��F� UT���Z ,<�TQ? b�y@�t�G?t�E� |�q>Q����[ ��Pa� RI��E� >SETUP2�_ \ �@=STD	p<TT������r��P�>RBACUbG] T��>R�d)�j�%C�E��0��IFI���0��i�{�4�PT�T��FLUI�D�^ Ђ gHPUR �gQ�"�r�a�4P�+ I�$��Sd�k?x��J�`CO�P��SVRT��N�x$�SHO* ��CAS�S��Qw%�pٴBG_%��3���<�FORC�B��^o�DATA��_�BKFU_�1�bb�2�apQn�b0��` |��wNAV	`�������$�S�Bu#$�VISI���2SCF	dSE�����V��-O�$&�BK�ἐ ��$PO��I���FMR2>��a �� �	��`#��&�8�PO� (�_���Ύ+IT_^�ۄ)M������DGCLFފDGDY�LD�����5Y&��Q$��M�됇Cb��{	 �T�FS�P�Dc �P��W�cK $E#X_WnW1%`]�Ԕ"X3�5��G�+�d ���S�WeUO�DEBU1G��-�GR��;@�U�BKU��O1nR� _ PO_ �)�����M��L�OOc>!SM� E��R�є�u _E �e � �TER�M`%fi%53,�'ORI�ae gi%�AGSM_�`>Re hi%�QV�(ii%UP>\Bj� -����e��w#� f��G��*ELTO�A�bF�FIG�2�a_����Ў$�$g$UFR�b$�1R0�օ� OT_7F�TA��p q3NST�`P�AT�q�0�2PTHIJ�ԀE�@�c3ART�P'5�Q�B΍aREL�:�aSHCFT�r�a�1�8_��QR��у�& � $�'�@i�
����s@bSSHI�0�Uy� �QAYLO�p�Oaq������1����pERV��XA��H��m7�`��2%�P�E3�P�RC<���ASYM�a�F�aWJ07����E���1�I��ׁUT�`Oa�5�F�5P�su@J��7FOR�`M ��G	RO!k]��5&�0�L0�THOL ;l� �s2T����OC�1!E�$OaP��qn���$�$����$��PR^��a�OU��3e��R��5e�X�1 �e$P�WR��IMe�BR�_�S�4�� �3�aU�D�ұ��Q�dm���$H�e!�`ADDR˶HR!G�2�a�a�aQ�R��[�n H��S����%��e3��e���e��SE��P��HS�MNu�o����Pªq��0O�L�s߰`ڵ�I A�CRO��&1��ND�_C�s��AfdK�R'OUP��R_�В� �Q1|�=�s���y %��y-��x���y���y�>�=A��Ҁ�AV#ED�w-��u,&s�p $_��P_D� ��'rPRM_�����HTTP_��H[�q (ÀOcBJ��b �$˶�LE~3�`��\�r G� ���ྰ_���TE#ԂS�PIC��K�RLPiHITCOU�!��L���PԂ�������PR��PSS�B�{�JQUERY�_FLAvs�@_W�EBSOC���HQW�#1��s�`<P�INCPUPr��O ���g�����d��t���O�T�IOLN.�t 8��R� ��$SL!$I�NPUT_U!$�`��Pw�֐SL.���u���2�.���C��B�0֐a�F_�AS=v�$L+ਇ+�A��bb41`�����Z@HYʷp����#qe�UOP:w `v�ϡ˶�¡�������"`PIC`����� �	�H�IP_sME��v�x Xv�cIP�`PrR�_N�p�d���Rʳp�ױ�QrSP �z�C��B�GPqL��M�Av�y3 l�@CTApB��AL TI�3UfP_ l۵�0PSڶBU_ ID� 
�L � `�0y���0z)����ϴ�NN�_ O���IRCA_CN�f� { �Ɖ6-�CYpEA���� ����IC�ǫ�tpR<�=QDAY_
��NTVA�����!�8�5����SCAj@��#CL�
����
����v�|5�VĬ2b�l�N_�PCV�n�
���w�})�T��S�����
���e���T� 2|C ��� �v�~�8�֣�ذLAB1��\_ ��UNIX���� ITY裪��ea��R� ��<)���R�_URL���$A;qEN ���s`vs�TeqT_U�� �iJ��X�M�$���E�ᒐR祪�� A��,���JH���FL�y��= 
���
�wUJR|U� �ƀAF�6G��K7��D>��$J7�s��J8B*�7���3�E�7���&�8\�)�APHI�Q4�y�DkJ�7J8R��L_K�E'�  �K�͐LMX� � �<U�XRi�����WATCH_VAZqxu@AំFIEL`�b�cy� ��:� � bu1VbwPCTX�j�n�LGE�߄� !��LG_SIZ΄�[8XZm�ZFDeIY p1!gXb ZW �S `�8�m��� ��b ��A�0_i0_�CMc3#�*'F Q1KW d(V(Bbpo pm�p� |Io�1 p�b pW RS��0 7 (C�LN�R��۠�DE6E�3����c�i���PL�#�DAU"%EA`q�͐�T8". GH�R���y�BOO�a��� C��F�IT0V�l$A0��RE���(GSCRX����D&�|ǒ�qMARGI4� Sp�,����T�"�y�	S��x�W�$y�$���JGM7MNCHLt�y�FN��6K@7�r�>9UFL87@L8F�WDL8HL�9STPL:VL8"�L8s L8�RS�9HOPh;��C�9D�3R��}P�'IU h�`4�'�5$ ��S2G09�pPOWG�:�%`�3,64��N9EX��TUI>5I� �ӌ������C3�C<0'�@,�o:��&�@�!Naq�vcANAy��Q�A�I]�gt7Ӝ�DCS����cRS�cRROXXO"dWS�ÂRoXS{X�(IGNp 
Ђ=10 ܰ�[TDEV�7LL ���y��C �	 8�Tr$f/蛒�Ĵ��3A�a�	 �W�萦�Oqs�S1
Je2Je3Ja��BSP�C � �ƋG`-T ��%��Q�T�r@�&�E�fST�R9 Y�Br�a �$E�fC�k�g��f	v�8lce�C � L���� � ��u�xs뀔�g�q��jt��!�#_ � [��w�#Ӡ �s� �MC�� =�ƀCLDP᠜�TRQLI ���y�tFL���rQ��s5�1D���w~�LD�u�t�uORG���1�?RESERV��M�Ⱥ�M�Œ�s��� � 	�u�5�t�u#SV��p��	1���}��RCLMC���M�_�ωА��;�MD�BGh�I����$�DEBUGMASP������U�$T8P���EF�d��pFR�QҤ� � ~K	HRS_RU4��bq��A��$EFR3EQ6u!$0YOVER�k��f��PU1EFI�!%Gq�� �7�
Y�z�ǐ \����E�$9U�`��?��
�SPSI`��	��CA ���ʲ�σUY�%��?( 	iaMIS�C�� d��aR5Q��	��TB� �c ���A��AX����𑧪�EXCESHg�!qd�M�Hᒅ�au���}qd�SC�`� � H�х�_������������pK�E��+�� &�B_^, FLICBtB� �QUIRE CMO�t�O���r�LdpMD� �p{!��5�b���$L�MND!��I����L� �D;
$INAU9T�!
$RSM���PN�b�C����PSTLH� 4nU�LOC�fRI"�v�eEX��ANG.R�.���ODA]��bq��� ���MF0 ����icr�@mu����$�SUPiuiaFX��IGG! � ���cs��#cs
F ct��ޒ�b5��`E��`�T�5�tC��g�TI���C`���M����� t�MD���) ��XP��ԁ��H��.���DIAa��Ӻ�W��!��0af���D@#)���pO�㥀��� -�CUp V	����.�֡O�!_��ᜃ ��p�c����	�� |�P|��0� ���P{�KEB��e-�$B��o�=pND2xւ����2_TXlt�XTRAXS����&��LO: ����}����C�.�&���RR2h���� -�!A�� ?d$CALI����GFQj�2F`RIN�bn�<$Rx�SWq0ۄ���ABC�ȇD_J��{�.���_�J3��
��1SPH, �.�P����3��(H�9p.�#J�34n���O�QIM�M�CSKP�zb7?SbJ+�M�Qb�y8����_AZ��/��EL�Q.ցOC�MP��N�� RTE�� �1�0 ����1��@ ZScMG�0����JG�p�SCLʠ��SPH�_�PM��f��.��u�RTER��n��Pk�_EP�q�`A0� �cM��DI�Q�23UdDF  쀐�LW�VEL��qINxr�@�_BALXP.��Y/�J�0�'$\�IN���B]�C�9%�".�
8!:6p_T� �F%a"�a�^$��k)�"p�DHʠ��\�9`�$Vw��_�A$�=��~�&A$���s�R6�]�H �$BEL� m���_ACCE� x	8�0IRC_��q�@�NT��c�$PSʠ�rL� ��M4�s9 .7��GP/6 ��9�7$3�73S2T�͡_Ga�"�0�1��8�n1_MG}�DD�1�~�FW�p��3�5�$32�8DEKPP�ABN[7ROgEE�2KaBO�p�Ka���1�$USE�_v�SP��CTR�TY4@� �� <qYNg�A�@�FR �ѢA!M:�N�=R�0O�v1�DINC(��B�4p���GY��ENC��L��.�K12��H0I�N�bIS28U��ON�T�%NT23_�~�fSLO�~�|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1���M�PERCH  �S��� �W���Sl� �R��l����E�0�0PAS2EeL�DP7��ONUЉZ�f�VTRK�RqAY"�?c� �aS2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gB�T�DUX �2S_BCKLSH_CS2 Fu:��V���C-�esR�oz�A�CLALM�JT@��`� �uCHK�e ����GLRTY@pн�8T��5���_��N�T_UM3��vC3�p�1Z���LMT���_LG��%���0�E *�K�=�)�@5F�@8 09�Nb��)hPC�Q)h�HТ��5�uCMC����0�7CN_��N����;SF�!iV �B��.W���S2/�Ĉ7CAT�~SH�Å� �4 V�q/q/V�T1���0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e�0�R� @B�_Wu�d��!a��#`��#`�I*h�Iv�I�#F��S��:��I�0VC00��֢1ܮ�0��JRKܬ!��<�KDBXMt�<�M��_DL�!_bGRV�g�`��#`��#A�H_p%�?��0��COS��� ��LN#���ߥŴ � ��=������꼰�b<�Z���VA�MYǱ�:ȧ��᯻[�THE{T0�UNK23�#؅��#ȰCB��CB�#Cz�AS�ѯ�0���#����SB�#��N��GTSkZAC�������&���$DU�phg6�j��E��%Q%a_��x�NE
hs1K�t�� y�A}Ŧկ׍������LPH����^U��S ߥ����������!�(�(Ʀ�V��V�غ ���V��V��V
�V��V&�V4�VB�H���������d�����H�
�H�H&�H4�H*B�O��O��Os���UO��O��O
�O�UO&�O4�O(�F����	���SPBALANCE_J��6LE��H_}�S�P>!۶^�^��PFULCb�q����K*1�UTOy_�p�uT1T2�	
22N�q2VP�M@�a� i�Z23	qTu`�O�1Q�INSE9G2�QREV�P�GQDIF�ep)1�lU�1��`OBK�qj�w2,�VP�qI�?LCHWAR4B�B�AB��u$ME�CH��J��A��vAX�aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ֯@�C1_ɒT �� x $W�EIGH�@w�$ȹ�\#��I�A�PIF�vA�0LAG�B��S��B:�BBIL�%O1D�`�Ps"ST0s"P:�pt � N�C!
L �P 
P2�Aɑ�  2��Tx&DEKBU�#L|0�"5�OMMY9C59N���$4w�$D|1 aq$0ېl� > �DO_:0AK!� �<_ �&� �q�A��B$�"� NJS�8_�P�@� �"O�p �� %�T7P?Q��TL4F0TICK,�#�T1N0%�3=pB�0N�P� u3�PR\p��A��5��5U0PR�OMP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a��@RU�COD�#F9U�@�&ID_�P�E�82B> G_SUFF�� �#�AXA�2DO�7/�5� �6GR�#��DC�D ��E��E-��DU4� u�_ H_FI�!�9GSORD�! R 236s�HR�A>N0$ZDT�E=!|� X5�4 *WL_NA�1�0�R�5DEF_I�X�RF �T�5�"�6�$�6�S�5�UFISm�#�m1|Ј�40c�3�T6�44􁆂�"D� ?rfd�#�D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D�S �D�U�D>b�B�c�E�S �Dd�B�&2v2a�C� ʑ�E�R�E�S�C9wwu�H�0P} d�0,a���F0W�h�u�c����TE�qY4�� �!LOMB�_�r�w0s"VIS���ITYs"AۑO>�#A_FRI��F~SI,a�n�R�0H7��07�3�#s"W�!W�Q��%�_���AEAS{#�B��|��x`WB8�45�55�6�|#ORMULA_�I���G�W� �h 
>75COEFF_O�1&)�$�1��Go�{#S� 52�CA� :?L3�!GR�m� � � �$�`�v2X�0TM��g���e�2�c��3E�RIT�d�T� � M �LL�Dp`S��g_SVkd��$�v�� �.���� � ޅ�SETU,cMEAG@�@Πt �!HRL �� � (�  0��l��l��aw�"�R�0�a�a}d]�Ad��B��Ay`Ga�x`��[Ѐk@RE�C[Qq��QSK_�A y�� P_!1_USER����p�*���VEL�� ��-�!��IzPBw�MT�1CFG����  �0]O�NOREJ �0l����[�� 4 �e���"�XYZ�<SB� 3����_7ERRK!� U ѐ�1�@c�Ȱ�!�>��B0BUFINDqX���p� MORy�7� H_ CUȱ�1���dAyQ?�I>Q'$ +�a������ \�G{�� � $SI�h��@�2	�VOv�q�- O�BJE| w�ADJ1UF2yĈ�AY�����D��OUKP���\�AMR=�Tp��-���X2DIR�����Xf�1  DYNHt�0�-�T� ��R���0� ���OPWO}R�� �,B0�SYSBU����SCOPo���z�Uy�bXP�`K���PA��q������OP�@U����}�"1��IMAG۱_ �п"3IM.���IN����~��RGOVRD"���	���P����  >PgplcC��L�`BŰ|?l�PMC_E�P�1N��Mr�12112�P"�SL| ���� �R OVSL:=S�rDEX\a`"��2�:�_"��� P#���P������2�C �P>���#�/_ZERl���:����� @��:��O&�@RIy��
[�g@�e���s�~�PL����  $FREEY�EU���Z���L����T�� A�TUSk�,1C_T�����B������p��Vc1��P��� Dc1�к���LQ����0MQ��ۡL�XE��x�5IP�W�` ��cUP��H`&aPX;@���43����PGY��g�$S�UB���q���J?MPWAIT~ ���LOW���1wē �CVF_A�0��RX�Z��CC �R$���28IGNR_P�L��DBTB� P�*a�BW@.t�UL�0-IG��!@I�OTNLN,�RB��b�N!@��PEE�D~ ��HADOW� ��t���E�����ܹ�PSPD��� L_ A�нP���	#CUNq � �RP F(�LYwPa����_PH_PK���b�?RETRIE��x���ҋRS D@FI���� ���V �$ 2}�d�DBGLV<?LOGSIZz�baKKTU���$D�n�_TXV�EM�!Cڡ)�� �-R�#�r>��CHECKz��(��L���ϰq)ҹL��NPA�`T(J"����*0P����
�AR�"�BC =S�a��O�@����ATTS�u䡳&� w�^a��3-#UX^�4�P9L�@Z�� $d��q?SWITCH�h�-W��AS��f�3�LLB��� /$BA�Dvc���BAMi��6I��F(@J5��N�UB6[F>
A_KNOWK3qB"�U��AD+Hc� �D��IPAYLOAq�9p�C_���Gr�*�GZ�CLqAj��P�LCL_6� !�4��BOA?�T7�
VFYCӐ�Jp��D
�I�HRՐ�G�T�B��6�J(�zQ_Jt�A �B�AND�����T�BQ}!��PL~@AL_ ��0� =�TAe��pC��D:�CE���J3�P�V�� T�PDCK�^�)b��COM�_AgLPH�ScBE<�߁�_�\ �X�x\�� � ���OD�_1�J2�DDM�A�R<�h�e�f�cQ�TWIA4�i5�i6��MOM(��c�c�c�c4�cV�B� AD�cv��cv�cPUBP�R �d<u�c<u�b}"�1����� L$PI $��pc��G�y��I*�yI�{I�{I�s�`@�A���v��v�J��b��a��HIG �3���0���5 �0�f�?�5N�5�SAMPD Ƣ�0�p���;@�S �� с6���1���� �� �`���`1�K�P��`�d�P�H��IN1� �P��8�T�/��:�z�xQ�z���GAMM&��S��$GET������D^d>�
$N�PIBR��I��$HI��_���1��E=��A�9�*�LW�W�N�9�{�*��Zb���QCdCH�K0�j�ݠnI_ ��M�JļRoh�Q ���sJ�-v��S {�$�X 1�N�}I�RCH_D�$RN���^�L�E��i�p�Zh8�ž�MSWFL/Mn�PSCR�75��� ��3�"Ķ�6��`���ع��f0jqSV��P'�������GRO�g�S_SaA=AH�=ńNO^`Ci�_d=��no�O �O�x�ʚ��p�B�u���cDO�A��!� ں�*�t�:�Z1f�;�x7����C �}Mmu� � �#YL�snQ ���  ���"��<s�	������nQ૰<3M_	Wl�����\p��(�o�MC��P���QA����hpM.�pr� ��!��$�yWM��ANGL�! �AM�6dK�=dK�DdK��TT7�Nk@��3�#J�PXC OEc�QZ��hp	nt� ���OM���ϑϣϵπ���`� c�Z0es^a_�2� |a�J��i ���c���cJ��j����8�jA� v�¥�{ �@{�P�1�PMON_QU��� � 860QCsOU��QTHxsHO��B HYS�03ESPBB UE- 3ºf0O�4�  c P��^�RUN_T�O��n��� �P�@��IND9E�#_PGRA���0���2��NE_NO���ITf��o INFO��a"��Θ���� =(*�SLEQ!�*0�*�I�OS��l4�� 460ENA�By� PTION��3��r��^GC]F�!� @60J�,�Q���R�d!���erPEDITN�� �� ��KAQj"� �E(�NU'�(AUTY�%CO�PYAQ�2,�qe�M��N< @+��PRU�Tm� C"N�OU��2$G��$erR�GADJ��u2X_��IX����&���&W�(P�(~��&9�� z
�N�P_CYCy�$RGNSc֜{�s�LGO£�NYQ_FREQSrAW@��X1�4�L�@��2P0�!�c@�"�CR1E��MàIF�q��NA��%�4_G>f�STATU~�f���MAIL��|CI<q�=LAST�1a�*4ELEMg� ���QrFEASI t;�ւΰ��B"�F�AF����I� ��O2`�E u�vBAB��PE� =�VA�FzQ��I��TqU[��R���S�FRMS_TRpC�Qc��C��Z�
�`�1�Ds�*4ns؆��	MB 2�  `���N�3V�R2WR*����шR^W�wj�DO�U�^�N�,2PR�`�h�1GRID���BARS!�T�YuZ�Op��+ |_�4!� �R�TO��d� � 9����POR�c\~vbSRV�0)"dfDI[�T�`;aNd�pXg
�Xg4Vi��Xg�6Vi7Vi8:afqF�ʒg�z $VALU�C0�3Dr�ad�� !pf��b�S�1-ȆAN/���b�1R�]11ATO�TAL����=sPW�E3I�QStREGENQzfr��X�H�]5	v( TR�CS�QqC_S3��wfp�V�!��r��BE�3�PGp0B�( sV_H�P�DA(��p�S_Yha���i6S��AR(��2� �"IG_CSE�3�pb�5_� ��tC_�V$CMP,l��DEp�G����IšZ~�X��R�aE�NHANC.� p Qr�2���GINT9`cq�F����MASK�3�@OVRMP �PD�1@-��W�QaХT�l�_RF�{�V�PSL)GP�g�9�j5��,�;pDpS���4���U����`�T9E���`���`k�ⵥJ^�Y�y3IL_�Mx4�s��p��TQ@( ���@����V.��C<�P_ �R�F�M�]�V1\�V1j�2�y�2j�3y�3j�4y�4j���p۲�������ܲIN�VIAB8�6�#��*�2&�U22�3&�32�4&�!42��6�I�SJ�  ��T $MC�_FK `� �LP>�J�х1pMj�Iу��zS ��1����KEEP_HNA�DD��!鴓@�C��0	��Q����
�O!�v ���p
�և.
�REM!�	�CqP�RF�]�b�U�4e	��HPWD  ��SBM���PCOLLAB*�p��/q�2IT/0��Q"{NO1�FCALp�܎���� , �FL|v�A$SYN����M��Ck��RpU_P_DLY��z�DELA9�Dq�2Y� AD(�'0�Q�SKIPO�� �4`� O��NT����c�P_� ��׾ �� cp���q�ٞ��o`�� |`�ډ`�ږ`�ڣ`����`��9�!�J2RT0  �lX�@TR3 H��1AH� �H����PRDCq���+ � R�R, 5���R�1��E��5TR�GE�_C��RFL�G"���W�5TSsPC�1UM_H��2TH2N}Q��;� 1� ��;��Q02 �� D� ˈ��@2_PC3W�S���1Y0_L10_Cw2���,��� � $ \� U@��V7������0��VU\�� ��� rd��C��+��*7��DZ Gs�RUVL1[�1h���;10]�_DS��7�����PK 11�� �lڰ����q��AT?��$�Q[7�� ���K 5T���HO�ME� *�c2h�n�����
�3h���!\3E `4h�hz����&0
`5h���	//(-/?/�6h�b/t/��/�/�/�/�7h���/�/??'?9? ���!8h�\?n?�?ؒ?�?�? ��FP�S����  @�Aa{p��]_�Ed� T=�nD4vnC�IO䑎II@`�O��_OP�E�C.r����POWE	��� X@�f���$$Cd�S�������A3�3� ��@�SI��G�P0�QI�RTUAL�O
QA�AVM_WRK �2 7U� 0  �5�Qn_zXk_�] �\	�P�]�_3�B8P��_�_�Ve�\ #m/o�Q5ojo|o�dHPsBS�� 1Y� <Xo �o�o�o�o#5G Yk}����� ����1�C�U�g� y���������ӏ��� 	��-�?�Q�c�u��� ������ϟ���� )�;�M�_�q�������й�˯ݯ�bC$�AXkLM�@���c7  d�IN�����PRE
�E��J�-�_UP��[��7QHPIOCNV_��� �	�Pr�U�S>��g�cIO)�Vw 1U[P $E`���Qս9lҿ8P?� � �����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y������� ��������	-? Qcu����� ��);M_ q������� //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo��o�o�o�o�o�m�L�ARMRECOV� a��-���L�MDG ���ɰ�LM_IF ���ை�� ��zv���%�6�?, 
 6�_���r漅�������̍$ w���׏��8�J�\��n����NGTOL�  a� 	 �A   ��ț�P�PINFO ={ <v����1��  I�3�a�"r P���t��������ί ���>�o����j� |�������Ŀֿ������0�B�PzPPL�ICATION �?����+�Hand�lingTool� �� 
V9.?30P/04ǐM�
88340����F0����202�ťʚϬ�7DF�3��M̎�None�M�FRAM� �6��Z�_ACoTIVE�b  s�  p�UTOMODz�A���m��CHGAPONL��� ��OUPL�ED 1ey� �������g�CU�REQ 1	e{ � T���	�p��w���#r����e��HN���{�HTT�HKY��$r��\ [�m����O�	�'�-� ?�Q�c�u��������� ����#);M _q����� �%7I[m ���/��� /!/3/E/W/i/{/�/ �/�/?�/�/�/?? /?A?S?e?w?�?�?�? O�?�?�?OO+O=O OOaOsO�O�O�O_�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ oo#o5oGoYoko}o �o�o�o�o�o�o 1CUgy�� �����	��-�`?�Q�c���1�TO���|�p�DO_CL�EAN��n��NMw  �� ��B�T�f�x���%�DS�PDRYR��m�H	I���@/����� ,�>�P�b�t�������8��ίj�MAXa�ۄ�������Xۄ����|��p�PLUGG�и܇�ӌ�PRC��B�� ��ׯF�OxK���ȔSEGF��K�������.������,�>�v���LAP ӟ澨�Ϥ϶����� �����"�4�F�X�j�>��TOTAL�7����USENUӰ��� ���ߖ�1�RGDISPMMC��e��C����@@Ȓ���Oѐ�����_�STRING 1�
��
�Mڥ�Sl�
A�_I�TEM1K�  n l�g�y�������� ����	��-�?�Q�c��u���������I�/O SIGNA�LE�Tryout ModeL��Inp��Sim�ulatedP��OutOV�ERRА = 1�00O�In c�yclP�Prog Abor�P���Statu�sN�	Heart�beatJ�MH� Faul��Aler�	�������*<N` ׃G�ׁY�c� ����////A/ S/e/w/�/�/�/�/�/8�/�/wWOR��G� -1�?U?g?y?�?�? �?�?�?�?�?	OO-O�?OQOcOuO�O�O�NPOE��@E;�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oop&o8oJo�BDEV�N u`�Obo�o�o�o�o�o �o,>Pbt��������PALT��E?� A�S�e�w��������� я�����+�=�O�pa�s����GRI� G뽑1������	�� -�?�Q�c�u������� ��ϯ����)�����R�a�՟;����� ����ѿ�����+� =�O�a�sυϗϩϻ�<��O�PREG�� y���-�?�Q�c�u߇� �߽߫����������)�;�M�_�q����$�ARG_-0D ?�	�������  	�$��	[��]���������SBN_CONFIG��� ��C�II_SAVE � ��)���TC�ELLSETUP� ��%  O�ME_IO����%?MOV_Hn������REPd�����U�TOBACKY����#�FRA:\�� ����)��'`l ��&�� 7"� �24/07/25� 10:26:54�����͓������+=Oas�Ƅ�� �����/1/C/ U/g/y/�//�/�/�/ �/�/	?�/-???Q?c?u?�?�?p���?�?�?��?�?	OO��OIN�I�Y�-���MESSAG9�GA)�|��RKODE_Ds�<��zHOw`�O���PAUS�@ !���� ,,		�����O�G�O__ #_%_7_q_[_�__�_��_�_�_�_�_%o����D�@TSK  ��M&,O��UPDT̀@EGd�`�FXW?ZD_ENBED��fSTADE��e���XIS�UNT �2��&�(�� 	\o��;&_ J�n�����d�METc�2LfE�� P�!��E��yS�CRDCFG 1��� �A�&�:�����ԏ�����Q=���H� Z�l�~�����	�Ɵ-� ���� �2�D��������GR�`�`�O��_UP_NA����s	��_EDC@�1n�� 
 ��%-BCKED�T-q����%�p���(��-��������������  ����2����t�� �d?���*�q���ϧ���3b�ҿ����΋�@��=�O���sϏ�4.� ��{����W���	����?ߏ�5��j�G�� �#������}�6��6��Z����Z� ���I��7��� ��&�λ�&m�������8^��*�� 	͇�9K�o��!9*�w��	�S���;��CR ����B/T//�/���w//��РNO_�DEL����GE_�UNUSE���I�GALLOW 1���   (�*SYSTEM�*)�	$SERV_GRǢ)�B0�@7REGK5$m3)��B0NUMp:�3�=�PMU� )�L�AY�p)�P�MPALD@�5CY'C10�.�>�0�>CULSU�?�=�2��AM3LOWDBO�XORIt5CUR�_D@�=PMCNmV�6D@10�>>�@T4DLI�`=O�_9	*PROGR�AJ4PG_M1I�>�OPAL�E_�UPB7_B>$�FLUI_RES�U�7p_z?�_�TMRY>h0�,�/�b�_�_ o o2oDoVohozo�o �o�o�o�o�o�o
 .@Rdv����������"LA�L_OUT �1;l���WD_AB�OR�0?d�ITR_RTN  �����g�NONST�OǠ�� 8CE?_RIA_I0���ۀ��ŀFCFG ��۔���_LIMY22�ګ �  �# 	i�J��<e�g�:�5�� 9��������
���u���PAQPGP 1�����Q�c��u�4�CK0����C1J��9��@���PC���CV��]��d��l­�s��P���C[�٤m��v���������� C�����-���?�ÂHE� ONFI�Pq�G��G_P�@1� �%�������ǿ�ٿ����G�KPA�USaA1�ۃ �2�W��Eσ�i� �Ϲϟ���������� #�I�/�m��eߣ���M��NFO 1v"��� �7���ߖ��� Dۊ��DH1�4 G ´-�?�ŀO��c�COL_LECT_�"�[�����EN�@��y�ܮ�k�NDE���"�3�"1234567890� �\1�� ��֕@�(��)M�r�\,L�^��� ]+������������C  2�Vhz� �����
c .@R�v��������� |����IO !����$���u/�/�/�/�C'TR�2"'-(�׀^)
��.R�#�R-�*W� 9_MOR�$� �;�l5� l9�?r?�?�?�?�;E2T��%S=,W�?@��@��C׀K)Dց
C�R�&u�XOWAWBVC�A�$��׀x׀�A"@Cz  Bʇ@C@�B8��AC�  @yB�׀�ց:d�43 <#�
�E��I�OT�C=AI��'GM?�C��(S=���Qd=AT�_DEFPROG �;%�/m_APINUSE�V�ۅ��TKEY_TBL�  s�ہ���	
��� !"�#$%&'()*�+,-./�:;�<=>?@ABC�DPGHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����Ga���͓��������������������������������������������������?������!�P�LCK�\���P�PS�TAn��T_AUT/O_DO��NFs�IND���n��R_3T1wT2N�����5ŀTRLCPL�ETE���z_S�CREEN ~�kcscÂ�U��MMENU ;1)O� <�[_ #�$��,�a���>�d� ��t���ӏ����	��� ��Q�(�:���^�p� ������̟�ܟ�;� �$�q�H�Z������� ���Ưد%����4� m�D�V���z���ٿ�� ¿�!���
�W�.�@� ��d�vϜ��ϬϾ�� ����A��*�P߉�`� r߿ߖߨ�������� =��&�s�J�\��� ���������'�,�p_MANUAL��EqDB
12�v�iDBG_ERRLIPs*�{h! 0�������g�NUMLIM�s:QOE�@�DBPXWORK 1+�{��>P�bt��-DBTB_�q ,��kC3!�VD!DB_A�WAYo�h!GC�P OB=��A�_CAL���o�k�Y�p�uO@`�_�� 1-
�+@
-k-6[l��_M+pIS�`��@"@�ONTImM�w�OD���&
�U;MOTN�END�_:REC�ORD 13�{� ��[CG�O� f!T/[K��/�/�/�/ _(�/�/f/?�/??Q? c?�/?�??�?,?�? �?OO�?;O�?_O�? �O�O�O�O(O�OLO_ pO%_7_I_[_�O_�O �__�_�_�_�_l_!o �_,o�_io{o�o�oo �o2o�oVo/A �oeP^�
�� �R���=��a� s��������*�ߏN� ��'���ԏ]�̏�� ������ɟ۟v���n� #���G�Y�k�}����TOLERENC��B�0� L���g�CSS_CNS�TCY 24	�t���.����� �0�>�P�b�x����� ����ο����(��:�äDEVICEw 25ӫ � �ϟϱ������������/�AߟģHND�GD 6ӫ� C�zT�.!ơLS 27t�S������������/�U�ŢPARAM 8Gb��A�Ք�RBT 2]:8�<����CkA� �·�  � �A���.SB����A�B�  ����������.�����  ����A�A�C����c�u����C�A�D���k�pz�A�A��HA�c��A�	�?( uL^p���A��Bt/�D��C���_ 	 A�=��ABffA�#33AҊ��g�A�A�Cf���a��A�J��7B�]��B��B�ffBᴠ�3�3C$.@R� (����A��� �
/��//)/;/ �/_/q/�/�/�/�/�/ �/�/<??%?r?I?[? m??�?�?�?�?�?&O 8O�PObOMO�OqO�O �O�O�O�O_�OO L_#_5_�_Y_k_�_�_ �_�_ o�_�_6ooo loCoUogo�o�o�o�o �o�o �o	h�O �w�����
� �.�	__I'�1_� q��������ˏݏ� ��%�r�I�[���� ������ǟٟ&���� \�3�E�W����ȯ�� �ׯ�"��F�1�j� E�s�����m������� ѿ�0���f�=�O� a�sυϗ��ϻ���� ����'�9�Kߘ�o� ������[����(�� L�7�p��m��� ��������$����� l�C�U���y������� ���� ��	V-? �cu����
 ��@+dO�s ��������*/ //`/7/I/[/m// �/�/�/�/?�/�/? !?3?E?�?i?{?�?�? �?�?�?�?�?FO�jO UOgO�O�O�O�O�O�O __�'O9OO=_O_ �_s_�_�_�_�_�_�_ �_oPo'o9o�o]ooo �o�o�o�o�o�o: #5��O��� �� ��$��H�Fz��$DCSS_S�LAVE ;����w���`�_4D  �w���AR_MEN/U <w� >�؏@���� �2�^rǏ�\�n�\���SHOW� 2=w� � fr[q����Ə��� ��,�>�D�b�t��� ����ҟϯ��� �)�P�M�_�q����� ����˿ݿ���:� 7�I�[ς�|Ϧ��ϵ� ��������$�!�3�E� l�fߐύߟ߱����� �����/�V�P�z� w����������� ��@�:�d�a�s��� ��������\���*� H�N�K]o��� �����28� GYk}���� ��"�1/C/U/ g/y/�/��/�/�/� �//?-???Q?c?u? �/�?�?�?�/�??O O)O;OMO_O�?�O�O �O�?�O�?�O__%_ 7_I_pOm__�_�O�_ �O�_�_�_o!o3oZ_ Woio{o�_�o�_�o�o �o�oDo-Se �o��o�������.�=�O���CFoG >������q��dMC:�\��L%04d.'CSV\��pc����m���A ՃCH݀�z�v�w�#��q���:�J�8�7����JP�j�)�́�p+�n�RC_O�UT ?z����a�_C_F�SI ?�� |���� �@�;�M�_������� ��Я˯ݯ���%� 7�`�[�m�������� ǿ�����8�3�E� Wπ�{ύϟ������� �����/�X�S�e� wߠߛ߭߿������� �0�+�=�O�x�s�� ������������ '�P�K�]�o������� ����������(#5 Gpk}���� � �HCU g������� � //-/?/h/c/u/ �/�/�/�/�/�/�/? ?@?;?M?_?�?�?�? �?�?�?�?�?OO%O 7O`O[OmOO�O�O�O �O�O�O�O_8_3_E_ W_�_{_�_�_�_�_�_ �_ooo/oXoSoeo wo�o�o�o�o�o�o�o 0+=Oxs� �������� '�P�K�]�o������� ����ۏ���(�#�5� G�p�k�}�������ş ן �����H�C�U� g���������دӯ� �� ��-�?�h�c�u� ��������Ͽ���� �@�;�M�_ψσϕ� ������������%� 7�`�[�m�ߨߣߵ� ���������8�3�E� W��{��������� �����/�X�S�e� w��������������� 0+=Oxs� ����� 'PK]o��� �����(/#/5/ G/p/k/}/�/�/�/�/ �/ ?�/??H?C?U3��$DCS_C_�FSO ?�����1 P [?U?�?�? �?�?�?O
OO.OWO ROdOvO�O�O�O�O�O �O�O_/_*_<_N_w_ r_�_�_�_�_�_�_o oo&oOoJo\ono�o �o�o�o�o�o�o�o' "4Foj|�� �������G� B�T�f���������׏ ҏ�����,�>�g� b�t���������Ο�� ���?�:�L�^����������ϯʯܯg?C/_RPI~>�?� ;�d�_�
�}?.�p���X�ݿj>SL�@�� �9�b�]�oρϪϥ� �����������:�5� G�Y߂�}ߏߡ����� �������1�Z�U� g�y���������� ��	�2�-�?�Q�z�u� ������������
 )RM_q�� �����*% 7Irm��� ��/�ϛ�,�/ W/�/{/�/�/�/�/�/ �/???/?X?S?e? w?�?�?�?�?�?�?�? O0O+O=OOOxOsO�O �O�O�O�O�O___ '_P_K_]_o_�_�_�_ �_�_�_�_�_(o#o5o Gopoko}o�o�o�o�o �o �oHCU g��������� ����NOCO�DE @������PRE_?CHK B��3��A 3��< �7��������� 	 <�����?# ۏ%�7��[�m�G�Y� ������ٟ�ş�!� ���W�i�C�����y� ïկˏ������A� S�-�_���c�u���ѿ �������=��)� sυ�_ϩϻϕ����� ���'�9���E�o�I� [ߥ߷ߑ��������� #����Y�k�E��� {����������� C�U��=�����w��� ������	����?Q +u�a���� ��);_q g�Y��S��� �%/�/[/m/G/�/ �/}/�/�/�/�/?!? �/E?W?1?c?�?�� �?�?o?�?O�?�?AO SO-OwO�OcO�O�O�O �O�O_�O+_=__I_ s_M___�_�_�_�_�_ �?�_'o9oo]oooIo �o�oo�o�o�o�o #�oGY3E�� {�����o� C�U��y���e����� ������	��-�?�� K�u�O�a�������� �͟��)��1�_�q� �}�������ݯ�ɯ �%���1�[�5�G��� ��}�ǿٿ����� ��E�W�1�{ύ�G�u� ���ϯ������/�A� �-�w߉�c߭߿ߙ� ��������+�=��a� s�M���ϑ����� ���'��3�]�7�I� ������������� ����GY3}�i �������� C/y�e�� �����-/?// c/u/O/�/�/�/�/�/ �/�/?)?�?_?q? K?�?�?�?�?�?�?�? O%O�?IO[O5OO�O kO}O�O�O�O�O_�O 3_E_;?-_{_�_'_�_ �_�_�_�_�_�_/oAo oeowoQo�o�o�o�o �o�o�o+7a W_i_��C��� ��'��K�]�7�i� ��m��ɏۏ����� ��G�!�3�}���i� ��ş������1� C��g�y�S�e����� �����ѯ�-��� c�u�O�������Ͽ� ןɿ�)�ÿM�_�9� kϕ�oρ����Ϸ�� ����I�#�5�ߑ� kߵ��ߡ������� 3�E���Q�{�U�g�� ����������/�	� �e�w�Q��������� ������+Oa �I������ �K]7� �m�����/ �5/G/!/k/}/se/ �/�/_/�/�/�/?1? ??g?y?S?�?�?�? �?�?�?�?O-OOQO cO=OoO�O�/�/�O�O {O�O_�O_M___9_ �_�_o_�_�_�_�_o o�_7oIo#oUooYo ko�o�o�o�o�o�O�o 3Ei{U�� ������/�	� S�e�?�Q�������я ㏽����O�a� ������q���͟���� ���9�K�%�W��� [�m���ɯ�����ٯ �5�+�=�k�}���� ���������տ�1� �=�g�A�Sϝϯω� ���Ͽ�������Q��c����$DCS_SGN CS������g��25-JUL-�24 10:30� EӘ� ����� X�S��������������Д�����Þ������  {�VE�RSION ���V4.2.�10�EFLOG�IC 1DS���  	�D���X�k�X�z�M�P�ROG_ENB � ��b��Л�U?LSE  ����M�_ACCLI�M��������WRSTJNT�����w�EMO���ѷ�L��INIOT EZ�O���OPT_SL ?�	S�1�
 	�R575�Ӆ�74*��6��7��5A��1��2��l���G�h�TO  t���.�H�V?�DEX��d����FPATHw A��A\4����HCP_CLNTID ?+�b� l������IAG_GRP� 2JS�_ ���[��D�  D��� D  B� w B�@ff�چ/B�@[��W��@�q��B��N�C�-BzBp@e`���mp3m7� 7890123�456�*�[�� � Ao�mA�j1AdA�]�
AW|�A�P�AJ-A�C/A;�A�4H���@�  �A��A�A3!_Ae�@@��B4��G ��t���
��uƨApffA�j�yAeK�A�_�AY��A�S� MC�AF��A@ �O�+/=/�O$O�c K�w(@�X�?8��@��y�/�/�/�/�/8��;d�2�5?@�~ff@x1'@�q��@kC�@�d�D@]��@Vv�6?H?Z?l?~?�8s�0l��@e�@^��@W�\)@O��@H��0?<@7K�@.V�?�?�?�?
O8_S@M00G<@�A��@<1@�5��@/l�@�(Ĝ@!�0�\NO`OrO�O�Ox'g� L_K�;_�_�__g_�_ �_�_�_o�_�_�_Yo�koIo�o�o+o�oX��"� 2�17A�@J>���R
q?�33�?Y��r��^J7'Ŭ2q63p�4�F>r��L�J@�p�Zr�
�=@�@�Qi�jq��@G Ah�@���@�T= c�<��]>*�H�>V>�3��>���J<����<�p�q�x���� �?� �C��  <(�U��; 4Vr�33��@,
���A@��?R�o D��mR�x���Q��t�� ��Z�Џ��؏�,��i�?�7N�>�(��>�@Z�=����J��G�v�G�@J�B�E�����a��@�ǐ@���@��@�Q�?L ��
�ŲI�P���&���'��@�K�����Ag�q�PC�  C���Cuy�
���ʯ ?����	�@�Գ�4���X��v���+��A�¿��� �����@�+�F���Iϗ�CT_CONFIG K�3���eg���STBF_TTS��
����"���t����{�MAU�����MSW_CF���L  K �O�CVIEW	�MI�U��㯛߭߿� ���������0�B� T�f�x�������� ������,�>�P�b� t�������������� ��(:L^p� �����  �6HZl~�������/��R%CB�N��!�� F/{/j/�/�/�/�/�/���SBL_FAULT O9*^�1GPMSK��7���TDIAG PԺ�U����q�UD1: 67�89012345 q2�q���%P�ϭ? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �a6�I'�
�?_�ƟTRECPJ?\:
 j4\_�7_[�?�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�O�O�_ _�UMP_OPTION��>q�TRB���9;uP�ME��.Y_TE�MP  È�g3B����p�A�pytUNI'��ŏq6��YN_BRK �Qt�_�EDITO�R q&qh�r_2PE�NT 1R9)  ,&�/0��d� [�`�J���n������� �ȏ��)�;�"�_� F�����|�����ݟğ ֟���7��F�m�T� ��x���ǯ���ү��!��E�,�i�P��pMGDI_STA�u�~��q�uNC_IN�FO 1SI��b�������Կⷮ�v��1TI� ��o(#��0�
0�d�o}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������Hu� � 2�D�R�j�R�x��� ������������,� >�P�b�t��������� ����Z��#5G a�k}����� ��1CUg y�������� 	//-/?/Yc/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?��?O%O7O Q/GOmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�? Ooo/o�_[Oeowo �o�o�o�o�o�o�o +=Oas�� ����_�_��'� 9�So]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�K�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�C�5�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� ������!�;�M�W� i�{���������� ����/�A�S�e�w� �������������� +E�Oas�� �����' 9K]o���� 1����/#/=G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?��?�? 	OO5/?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�?�_�_oo-O#o Io[omoo�o�o�o�o �o�o�o!3EW i{����_�_� ���7oA�S�e�w� ��������я���� �+�=�O�a�s����� ����ߟ���/� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������͟׿ ����'�1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߫�ſ�������� �;�M�_�q���� ����������%�7� I�[�m�������߯� �������)�3EW i{������ �/ASew ���������/ !+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?/� �?�?�?�?/#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�?�_�_�_�_ Oo-o?oQocouo�o �o�o�o�o�o�o );M_q���_ ����	o�%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�����ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߩ������� �����1�C�U�g� y������������ 	��-�?�Q�c�u��� �߫����������� );M_q��� ����%7 I[m����� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? ���?�?�?�?�O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�?�?�_�_ �_�_�?�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y�_�����_� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q��y��� ��˟�۟��%�7� I�[�m��������ǯ ٯ����!�3�E�W��i��� �$ENE�TMODE 1U��� + ���������»��RROR_P�ROG %��%������TABL/E  ���Q��c�uσ��SEV_�NUM ��  �������_�AUTO_ENB�  ̵��ݴ_N�O�� V�������  *����J����������+����(�:���FLTR����HIS�Ð������_ALM 1W.�� ����̍�+;����������0�?�_����  ���²u꒰TC�P_VER !�!��@�$EXTLOG_REQv�s�����SIZ����STK��������TOL  ���Dz~��A ��_BWDU�*�Z��V�ǲ?�DID� X�Z�����[�STEPl�~���>��OP_DO����FACTORY_�TUNv�d��DR_GRP 1Y��`�d 	p�.° ��*u����RHB ��2� ��� �e9 ���bt� o��������J5nY@��SQAYM�@I�Cm@�`�u
 E�����u ȸo��_/�(/(oB�  F!A��w�33R"�33-/@UUTn*@� �/ȷ>u.�>*?��<��ǆ-��F@ �"�5W��%�-J��NJk��I'PKHu���IP�sF!����-?�?�/9��<9�8�96C'6<,5���/�_?��FEATUROE Z�V�Ʊ�Handl�ingTool ��5��Engl�ish Dict�ionary�74�D St�0ard��6�5Analog� I/O�7�7gle Shift O�uto Soft�ware Upd�ate%Imati�c Backup��9SAground� Edit�0�7C_amera�0F�?�CnrRndIm�XC�Lommon �calib UI�C�FnqA�@Monoitor�Ktr�0?Reliab@�8�DHCP�IZat�a Acquis��CYiagnos�OA�1[ocume�nt Viewe��BWual Ch�eck Safe�ty�A�6hanc�ed�F�:�UsnPF�r�@�7xt. D7IO �@fiRT�Wwend�PErr�@QLQR�]�Ws�Yr�0��P E�:FCTN_ Menu�Pv S�8gTP In'`f�acNe�5GigE�`nrej@p Mas_k Exc�Pg�W�HT^`Proxy� SvoT�figh�-Spe�PSki�D�eJP�Pmmun�icN@ons�hu�rE`'`_�1abconnect 2x�ncr``struH�2z>peeQPJQU��4KAREL C�md. L�`ua��husRun-Ti��PEnvkx(`el� +R@sP@S/W��7License��Sn\�PBook(System)�:MACROs,�b?/Offse@�uaH�P8@_�pMR�@��BP^MechSt�op�at.p6R�ui�RKj�x�P�0P@)��od@witchȘ�>�EQ.���Op�tmЏ>��`fil�n\=�gw�uult�i-T�`tC�9PC�M funHwF�o�3T�R?�f�Regi��pr�`I�rigPF�V����0Num S�elb����P Ad�ju�`���J�t�atu��
�iZ�5R�DM Robot>�0scove�1F��ea7��PFreq� Anly�gRe�m`��Qn�7F�R�S�ervo�P���8S�NPX b�rNSN^`ClifQɮB�Libr�3鯢0 �q�����o�ptE`sGsag?��4�� -C���;��/I_mB�M�ILIBk�E�P OFirm6BU�PEc�Acck@sKTPT9X_C�eln����F��1�V�orqu>@imula�A�A�u��Pa�qU�j@t�Ã&�`ev.B��.@riP޿USB port �@�iP�PagP��R �EVNT�ϗ�nexcept�P��t�X�ſX�]VC�Ar�b�bf�V2PҦ�$�����SܠSCصV�S�GEk�a�UI�;Web Pl!��ާ���Խ`�TeQfZD?T Appl�d�:x�ƺ� �GridV�play�R�WD4�R
�.�:n�EQ+��r�-10iA/7L�*��1Graphi�c���5dv�SDC�SJ�ck�q�5la�rm Cause�/��ed�8Asc�ii�a��Load�nP�Upl,�Ol�0�AGu�6N�`���yFyc@�r�����P�V��Jo��m� c��R���c���m�./������Q�2*u:eRA`J��P�ٶ4eqinL�����8NRT��9O}n�0e Hel�H�J�`oI�allet�iz?�H�����_�t�r�[ROS Eth�q��T@e�ׅ�!��n�%�2D�tPkgp&Upg~��(2DV-�3D� Tri-jQEA�ưDef.qEBa)pdei��� �b�ImπF�f��n�sp.q=�464M?B DRAMZ,#�FRO5/@ell��<�Mshf!r/�'c�%3@pLƖ,ty�@s˒xG��m��. [�� ��BU���Q�B�=mai�P߫�]hQ����@q6wlu��H��^`�xR�?eL� Sup������0�P�`cr��@�R���b�x���pr1uest�Crt~QQ��ߋL!��4O��q$�K��l� Bui7�n��A'PLCOO�EVl%��sCGU�OCRG�Ob��DR��O
TLS_&��BU/_��K�qN_&d�TA�OxVB�_�Wp�ܑZ���_TCB�_ �V�_�W���WF+o�V��O�W._�W�ņoTE�H�o�f�O�gt�oT	Ej�xVF�_w�_xV�GoTwBTw~oxVH�xVIA��v�xVLN�yUMz�boH�f_xVN�xVP�H��^xVR&xVS��܇ʏ��W��v���gVGF:�L�P2_�h��h�V�h��_g�D���h�FFoh��g�R�D�� TUT��0�1:�L�2V�L�TB�GG��v�rain�UI��
%HMI���pon��m��f�"�F�&K�AREL9� �TPj��<5�
"E�<�N� {�r���������̿޿ ���A�8�J�w�n� �ϭϤ϶�������� �=�4�F�s�j�|ߩ� �߲���������9� 0�B�o�f�x���� ���������5�,�>� k�b�t����������� ����1(:g^ p�������  -$6cZl� �������)/  /2/_/V/h/�/�/�/ �/�/�/�/�/%??.? [?R?d?�?�?�?�?�? �?�?�?!OO*OWONO `O�O�O�O�O�O�O�O �O__&_S_J_\_�_ �_�_�_�_�_�_�_o o"oOoFoXo�o|o�o �o�o�o�o�o KBT�x��� ������G�>� P�}�t�������׏Ώ �����C�:�L�y� p�������ӟʟܟ	�  ��?�6�H�u�l�~� ����ϯƯد���� ;�2�D�q�h�z����� ˿¿Կ���
�7�.� @�m�d�vψϚ��Ͼ� �������3�*�<�i� `�r߄ߖ��ߺ����� ���/�&�8�e�\�n� ������������� +�"�4�a�X�j�|��� ������������' 0]Tfx��� ����#,Y Pbt����� ��//(/U/L/^/ p/�/�/�/�/�/�/�/ ??$?Q?H?Z?l?~? �?�?�?�?�?�?OO  OMODOVOhOzO�O�O �O�O�O�O_
__I_ @_R_d_v_�_�_�_�_ �_�_oooEo<oNo `oro�o�o�o�o�o�o A8J\n �������� �=�4�F�X�j����� ��͏ď֏����9� 0�B�T�f�������ɟ ��ҟ�����5�,�>� P�b�������ů��ί ����1�(�:�L�^����   �H552}���21n��R78��50���J614��ATU]PͶ545͸6���VCAM��CRIn�UIFͷ28	ƷNRE��52��R�63��SCH��DwOCV]�CSU���869ͷ0ضEI�OC9�4��R69���ESET���J�7��R68��MA{SK��PRXY!�]7��OCO��3�h����̸3�J6˸�53��H2�LCH^��OPLG�0֯MHCR��S{�MkCS�0��55ض�MDSW���OP��MPR�M�@�0n̶PCM �R0���ض��@�51�5u1<�0�PRS�ǻ69�FRD�FwREQ��MCN��{93̶SNBAE�^3�SHLB��M��tM���2̶HTC��TMIL����TP�A��TPTX��EL��Ѐ�8������wJ95,�TUT׻95�UEV��U�EC��UFR�V�CC��O��VIP��CSC,�CSGt8�r�I��WEB�7HTT�R6C�N��CGIG��IP�GS)RC�DG��H77��6ضR�85��R66�Ru7��R:�R530�K680�2�q�J��*H�6<�6,�RJح�j0�4�6o64\��5�NVD��R6��R84Tg�����8�90\���J9&3�91� 7+����,�D0oF�CL9I���CMS�� n�STY��TO䶴q���7�NN�O�RS��J% ��j�O]L(END��L���Sf(FVR��V3�D���PBV,�A�PL��APV�C�CG�CCR|�C�D��CDL@CS�Bt�CSK��CT�CTBL9��U0,(�C��y0L8C��TC� �y0�'TC(7TC���CTE\��07T�Eh��0��TFd8FJ,(GL8GI�8H�8�I��E@�87�CTM�,(M�8M@8N�8P�HHPL8Rd8(TSrd8W�I@VGF�GP2��P2���@�H�{7VPD�HF �V�PSGVPR�&VT���YP��VTB7Vs�IH��VI aH'VK��V���_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U?�g?y?�9  H55hT�1�1[Un�3R78�<50�9�J614�9ATU\�T�4545�<6�9�VCA�D�3CRIf,KUI8T�528-J�NRE�:52JR�63�;SCH�9D�OCV�JCU�48�69�;0�:EIOt�TsE4�:R69J�ESET�;KJ7�KR68�JMAS�K�9PRXYML7.�:OCO\3�<�J�)P�<3|ZJ6�<5u3�JH�\LCH\Z�OPLG�;0�ZM�HCR]ZSkMC�S�<0,[55�:MgDSW}k�[OP�[GMPR�Z�@�\0�:7PCMLJR0�k)P��:)`�[51K51�|0JPRS[6�9|ZFRD<JFR�EQ�:MCN�:9=3�:SNBA}K�[/SHLB�zM�{�@�ll2�:HTC�:T�MIL�<�JTPA��JTPTX�EL��z)`�K8�;�0�JJ�95\JTUT�[9�5|ZUEVZUE�C\ZUFR<JVCuC��O<jVIP,�wCSC\�CSGlJ��@I�9WEB�:H�TT�:R6{L��C�G{�IG[�IPGmS��RC,�DG�[�H77�<6�:R8�5�JR66JR7�[R|R53{6%8|2�Z�@Jml,|6|6\JR�\	P|�4L�6�64��5n�kNVDZR6+k�R84<���IP,�8f��90���KJ9�\91��̫7[KIP\J�D0�F��CLI�lKCMS�J9��:7STY,�TO�:�@��K7�LNN|ZOR�S<jJ��MZZ|OL�K�END�:L�S��FVR�JV3D�,�KKPBV\�AP�L�JAPV�ZCC�G�:CCRjCD��CDL̚CSBn�JCSK�jCTK��CTB��\���\�Ch�z���CL�TCLJl�l�TC��TCZ�CTE�J��|�TEX�J��<�TF��F\̥G��G��l�Hl�Ip�z)�l�k�CTM\�UM\�M��Nl�P,�eP��R��;�TS�ܹW��̚VGF��P2��P2�z ��VPDFLJVPn;�VPR��VT�;\� �JVTB��V�K�IH�VِM�<�VK,�V{��8#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew ������� +=Oas�� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G?�Y?k?}?�5�0�STD�4LANG�4�9�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~��������� �2�D�V�RB=T�6OPTNm�� ������Ǐُ���� !�3�E�W�i�{�����8��ß�5DPN�4� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳ڈ8�� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s���������pͯ߯��  ���*�<�N�`�r���9�9���$FEAT�_ADD ?	��������  	��ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu�����DEMO Z��?   ���} ��'��0�]�T�f� �������������� #��,�Y�P�b����� ������������ (�U�L�^��������� ���ܯ���$�Q� H�Z���~�������� ؿ��� �M�D�V� ��zόϦϰ������� �
��I�@�R��v� �ߢ߬��������� �E�<�N�{�r��� �����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo~o �o�o�o�o�o�o�o! *WN`z�� �������&� S�J�\�v��������� �ڏ���"�O�F� X�r�|�������ߟ֟ ����K�B�T�n� x�������ۯү�� ��G�>�P�j�t��� ����׿ο���� C�:�L�f�pϝϔϦ� ������	� ��?�6� H�b�lߙߐߢ����� ������;�2�D�^� h����������� ��
�7�.�@�Z�d��� �������������� 3*<V`��� �����/& 8R\����� ����+/"/4/N/ X/�/|/�/�/�/�/�/ �/�/'??0?J?T?�? x?�?�?�?�?�?�?�? #OO,OFOPO}OtO�O �O�O�O�O�O�O__ (_B_L_y_p_�_�_�_ �_�_�_�_oo$o>o Houolo~o�o�o�o�o �o�o :Dq hz������ �
��6�@�m�d�v� ������ُЏ��� �2�<�i�`�r����� ��՟̟ޟ���.� 8�e�\�n�������ѯ ȯگ����*�4�a� X�j�������ͿĿֿ ����&�0�]�T�f� �ϊϜ����������� �"�,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/
??A? 8?J?w?n?�?�?�?�? �?�?�?OO=O4OFO sOjO|O�O�O�O�O�O �O__9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿����&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t����������   ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�����y  �x�q��� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p��P����q�p�x ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p���������������$F�EAT_DEMO�IN  ��� �����IND�EX���I�LECOMP �[���B���8 SETU�P2 \B~L�  N w�5_AP2BCK� 1]B	  #�)����%����E �	���5 �Y�f��B ��x/�1/C/� g/��/�/,/�/P/�/ t/�/?�/??�/c?u? ?�?(?�?�?^?�?�? O)O�?MO�?qO O~O �O6O�OZO�O_�O%_ �OI_[_�O__�_�_ D_�_h_�_�_
o3o�_ Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0����ׯQ	� P� 2>� *.VRޯ(���*+�Q���W�{��e��PC������OFR6:��ؾg�����T   �2�����\� ��d�*.F��ϕ�	ó����qo�ߓ�STM� 9���ư%�d��ψ���HU߻�Jש�f�x���GIF�A�L��-����ߑ��JPG ����Lձ�n�����#JS�H�����6����%
JavaS�criptt���C�Se���Kֹ�v� %�Cascadi�ng Style Sheets���j�
ARGNAMOE.DT'��OЁ\;��[�k|(>k DISP*rU�Oп��� �
�TPEINS.X3ML/�:\C�cCustom Toolbar���	PASSWOR�D���FRS:�\�� %Pa�ssword Config/c�Q/ �J/�/���/:/�/�/ p/?�/)?;?�/_?�/ �??$?�?H?�?l?�? O�?7O�?[OmO�?�O  O�O�OVO�OzO_�O �OE_�Oi_�Ob_�_._ �_R_�_�_�_o�_Ao So�_woo�o*o<o�o `o�o�o�o+�oO�o s��8��n ��'���]���� �z���F�ۏj���� ��5�ďY�k������ ��B�T��x����� C�ҟg�������,��� P���������?�ί �u����(���Ͽ^� 󿂿�)ϸ�M�ܿq� ��ϧ�6���Z�l�� ��%ߴ��[����� �ߵ�D���h����� 3���W����ߍ��� @����v����/�A� ��e������*���N� ��r�����=��6 s�&��\� �'�K�o� �4�X��� #/�G/Y/�}//�/ �/B/�/f/�/�/�/1? �/U?�/N?�??�?>? �?�?t?	O�?-O?O�?�cO�?�OO(O�O�F��$FILE_DG�BCK 1]����@��� < �)
S�UMMARY.DyG�OsLMD:�O�;_@Diag� Summary�<_IJ
CONSLOG1__&Q_�_NQ�Console� log�_HK	T�PACCN�_o%�o?oJUTP A�ccountin��_IJFR6:I�PKDMP.ZI	PsowH
�o�oKU[`�Exceptio�n�oyk'PMEMCHECK5o�_*_K��QMemory� DataL�F�/l�)6qRIP�E�_$6�Zs%��q Packe�t L�_�DL�$y�	r�qSTAT����S� %~�rStatusT��	FTP���:����Vw�Qmmen�t TBD؏� �>I)ETHERNE���
q�[��NQEthern��p�Pfigura��oODDCSVRAF̏��ďݟd���� verify �all��{D�.���DIFF՟��͟xb��s��diffd���
q��CHG01 Y�@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ��VTRNDIAG.LS�̿޿s�^q=3� Ope���q� SQnostic�EWh�)VD;EV7�DATt�Q�xc�u�g�Vis��?Device�Ϫ�IMG7ºo����y�z�s�Imag�n��UP��ES��~T�FRS:\��� �OQUpdates List ��IJg�FLEXEVENQ�X�j߃�f��F� UIF E�v���B,�s��)
PSRBWLOD.CM��sL�������PPS_RO�BOWEL��GL�o�GRAPHIC�S4Dy�b�t���%4D Gra�phics Fi�leu��AOɿ��rGIG���u�
>YvGigE�ة�~�BN�? )��HADOW������\sShadow Chang���vbQRCMERR�n�\s�� CFG Er�ror�tail�� MA��C?MSGLIB� �"^o� ���T�)�ZD�����/XwZD�6 ad�HPNOTI���
/�/Zu�Notific8��H/��AGUO�/ yO?�O'?P?OOt?? �?�?9?�?]?�?O�? (O�?LO^O�?�OO�O 5O�O�OkO _�O$_6_ �OZ_�O~_�__�_C_ �_�_y_o�_2o�_?o ho�_�oo�o�oQo�o uo
�o@�odv �)�M��� ��<�N��r���� ��7�̏[������&� ��J�ُW������3� ȟڟi�����"�4�ß X��|������A�֯ e�����0���T�f� ���������O��s� �ϩ�>�Ϳb��o� ��'ϼ�K����ρ�� ��:�L���p��ϔߦ� 5���Y���}���$�� H���l�~���1��� ��g���� �2���V� ��z�	�����?���c� ��
��.��Rd�� ���M�q �<�`��� %�I��/� 8/J/�n/��/!/�/ �/W/�/{/?"?�/F? �/j?|??�?/?�?�?��$FILE_F�RSPRT  ����0�����8MDON�LY 1]�5�0� 
 �)M�D:_VDAEX?TP.ZZZ�?�?�_OnK6%N�O Back f�ile 9O�4S�6Pe?�OOO�O�?�O __?>_�Ob_t__�_ '_�_�_]_�_�_o(o �_Lo�_po�_}o�o5o �oYo�o �o$�oH Z�o~��C� g��	�2��V�� z������?�ԏ�u��
���.�@��4VIS�BCKHA&C*�.VDA�����F�R:\Z�ION\�DATA\v�����Vision VD�B��ŏ��� '�5��Y��j���� ��B�ׯ�x����1� ��үg�������X��� P��t���Ϫ�?�ο c�u�ϙ�(Ͻ�L�^� �ς��)���M���q�  ߂ߧ�6���Z���� ��%��I�������:�LUI_CONF�IG ^�5|m��� $ h� �3��������/�A�D$ |xq�s��� ��������a���  $6��Gl~�� �K��� 2 �Vhz���G ���
//./�R/ d/v/�/�/�/C/�/�/ �/??*?�/N?`?r? �?�?�???�?�?�?O O&O�?JO\OnO�O�O )O�O�O�O�O�O_�O 4_F_X_j_|_�_%_�_ �_�_�_�_o�_0oBo Tofoxo�o!o�o�o�o �o�o�o,>Pb t������ ��(�:�L�^�p��� �����ʏ܏��� $�6�H�Z�l������ ��Ɵ؟ꟁ�� �2� D�V�h���������¯ ԯ�}�
��.�@�R� d�����������п� y���*�<�N�`��� �ϖϨϺ�����u�� �&�8�J���[߀ߒ� �߶���_������"� 4�F���j�|���� ��[�������0�B� ��f�x���������W� ����,>��b t����O���(:�  �xFS�$FL�UI_DATA �_������uRESULT 2`��� �T��b����/"/ 4/F/X/j/|/�/�/� ��/�/�/�/?"?4? F?X?j?|?�?�?�?�=}?� 0�� ��?�;��O-O?O QOcOuO�O�O�O�O�O �O�O�#
O_/_A_S_ e_w_�_�_�_�_�_�_�_���?g�?;o �?boto�o�o�o�o�o �o�o(:L]o p�������  ��$�6�H�oi�+o ��Oo��Ə؏����  �2�D�V�h�z����� ]ԟ���
��.� @�R�d�v�����Y��� }�߯�����*�<�N� `�r���������̿޿ 𿯟�&�8�J�\�n� �ϒϤ϶������ϫ� �ϯ1�C��j�|ߎ� �߲����������� 0�B��f�x���� ����������,�>� ��G�!�k���W߼��� ����(:L^ p��S����  $6HZl~ �O���s�����/  /2/D/V/h/z/�/�/ �/�/�/�/�
??.? @?R?d?v?�?�?�?�? �?�?����9O� `OrO�O�O�O�O�O�O �O__&_8_�/\_n_ �_�_�_�_�_�_�_�_ o"o4oFoOO)O�o MO�o�o�o�o�o 0BTfx�I_� ������,�>� P�b�t�����Woio{o ݏ�o��(�:�L�^� p���������ʟܟ� ��$�6�H�Z�l�~� ������Ưدꯩ�� ͏/��V�h�z����� ��¿Կ���
��.� @�Q�d�vψϚϬϾ� ��������*�<��� ]����C��ߺ����� ����&�8�J�\�n� ���Q϶��������� �"�4�F�X�j�|��� M߯�q����ߗ� 0BTfx��� �����,> Pbt����� ���/��%/7/�^/ p/�/�/�/�/�/�/�/  ??$?6?�Z?l?~? �?�?�?�?�?�?�?O  O2O�;//_O�OK/ �O�O�O�O�O
__._ @_R_d_v_�_G?�_�_ �_�_�_oo*o<oNo `oro�oCO�OgO�o�o �O&8J\n �������_� �"�4�F�X�j�|��� ����ď֏�o�o�o�o -��oT�f�x������� ��ҟ�����,�� P�b�t���������ί ����(�:���� ��A�����ʿܿ�  ��$�6�H�Z�l�~� =��ϴ����������  �2�D�V�h�zߌ�K� ]�o��ߓ���
��.� @�R�d�v����� �������*�<�N� `�r������������� ������#��J\n �������� "4EXj|� ������// 0/��Q/u/7�/�/ �/�/�/�/??,?>? P?b?t?�?E�?�?�? �?�?OO(O:OLO^O pO�OA/�Oe/�O�/�O  __$_6_H_Z_l_~_ �_�_�_�_�_�?�_o  o2oDoVohozo�o�o �o�o�o�O�o�O+ �_Rdv���� �����*��_N� `�r���������̏ޏ ����&��o/	S� }�?����ȟڟ��� �"�4�F�X�j�|�;� ����į֯����� 0�B�T�f�x�7���[� ��Ͽ������,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸��߉��� ����!��H�Z�l�~� �������������  ���D�V�h�z����� ����������
. �����s5��� ���*<N `r1������ �//&/8/J/\/n/ �/?Qc�/��/�/ ?"?4?F?X?j?|?�? �?�?�?��?�?OO 0OBOTOfOxO�O�O�O �O�O�/�O�/_�/>_ P_b_t_�_�_�_�_�_ �_�_oo(o9_Lo^o po�o�o�o�o�o�o�o  $�OE_i+_ ��������  �2�D�V�h�z�9o�� ��ԏ���
��.� @�R�d�v�5��Y�� }�����*�<�N� `�r���������̯�� ���&�8�J�\�n� ��������ȿ��鿫� ���F�X�j�|ώ� �ϲ����������� ݯB�T�f�xߊߜ߮� ����������ٿ#� ��G�q�3Ϙ����� ������(�:�L�^� p�/ߔ�����������  $6HZl+� u�O������  2DVhz�� ������
//./ @/R/d/v/�/�/�/�/ }���?�<?N? `?r?�?�?�?�?�?�? �?OO�8OJO\OnO �O�O�O�O�O�O�O�O _"_�/�/?g_)?�_ �_�_�_�_�_�_oo 0oBoTofo%O�o�o�o �o�o�o�o,> Pbt3_E_W_�{_ ����(�:�L�^� p���������woɏ�  ��$�6�H�Z�l�~� ������Ɵ�矩� �2�D�V�h�z����� ��¯ԯ���
��-� @�R�d�v��������� п�����ן9��� ]���ϖϨϺ����� ����&�8�J�\�n� -��ߤ߶��������� �"�4�F�X�j�)ϋ� Mϯ�q�s������� 0�B�T�f�x������� �������,> Pbt����{� �����:L^ p�������  //��6/H/Z/l/~/ �/�/�/�/�/�/�/? ��;?e?'�?�? �?�?�?�?�?
OO.O @OROdO#/�O�O�O�O �O�O�O__*_<_N_ `_?i?C?�_�_y?�_ �_oo&o8oJo\ono �o�o�o�ouO�o�o�o "4FXj|� ��q_�_�_�_	��_ 0�B�T�f�x������� ��ҏ�����o,�>� P�b�t���������Ο ��������[� ���������ʯܯ�  ��$�6�H�Z��~� ������ƿؿ����  �2�D�V�h�'�9�K� ��o�������
��.� @�R�d�v߈ߚ߬�k� ��������*�<�N� `�r�����y��� ������&�8�J�\�n� ���������������� !�4FXj|� �������� -��Q�x��� ����//,/>/ P/b/!�/�/�/�/�/ �/�/??(?:?L?^? ?A�?eg?�?�?  OO$O6OHOZOlO~O �O�O�Os/�O�O�O_  _2_D_V_h_z_�_�_ �_o?�_�?�_o�O.o @oRodovo�o�o�o�o �o�o�o�O*<N `r������ ���_o�_/�Y�o ��������ȏڏ��� �"�4�F�X�|��� ����ğ֟����� 0�B�T��]�7����� m�ү�����,�>� P�b�t�������i�ο ����(�:�L�^� pςϔϦ�e�w����� �Ͽ�$�6�H�Z�l�~� �ߢߴ��������߻�  �2�D�V�h�z��� ����������
����� ��O��v��������� ������*<N �r������ �&8J\� -�?��c����� /"/4/F/X/j/|/�/ �/_�/�/�/�/?? 0?B?T?f?x?�?�?�? m�?��?�O,O>O PObOtO�O�O�O�O�O �O�O_O(_:_L_^_ p_�_�_�_�_�_�_�_  o�?!o�?EoOlo~o �o�o�o�o�o�o�o  2DV_z�� �����
��.� @�R�os�5o��Yo[� Џ����*�<�N� `�r�������g̟ޟ ���&�8�J�\�n� ������c�ů����� ��"�4�F�X�j�|��� ����Ŀֿ������ 0�B�T�f�xϊϜϮ� �������ϵ���ٯ#� M��t߆ߘߪ߼��� ������(�:�L�� p�����������  ��$�6�H��Q�+� u���a���������  2DVhz�� ]�����
. @Rdv��Y�k� }������/*/</N/ `/r/�/�/�/�/�/�/ �/�?&?8?J?\?n? �?�?�?�?�?�?�?�? ���CO/jO|O�O �O�O�O�O�O�O__ 0_B_?f_x_�_�_�_ �_�_�_�_oo,o>o PoO!O3O�oWO�o�o �o�o(:L^ p��S_����  ��$�6�H�Z�l�~� ����aoÏ�o珩o�  �2�D�V�h�z����� ��ԟ���	��.� @�R�d�v��������� Я������׏9��� `�r���������̿޿ ���&�8�J�	�n� �ϒϤ϶��������� �"�4�F��g�)��� M�O����������� 0�B�T�f�x���[� ����������,�>� P�b�t�����W߹�{� ������(:L^ p������� ��$6HZl~ ���������� ��/A/h/z/�/�/ �/�/�/�/�/
??.? @?�d?v?�?�?�?�? �?�?�?OO*O<O� E//iO�OU/�O�O�O �O__&_8_J_\_n_ �_�_Q?�_�_�_�_�_ o"o4oFoXojo|o�o MO_OqO�O�o�O 0BTfx��� ����_��,�>� P�b�t���������Ώ ���o�o�o7��o^� p���������ʟܟ�  ��$�6��Z�l�~� ������Ưد����  �2�D���'���K� ��¿Կ���
��.� @�R�d�vψ�G��Ͼ� ��������*�<�N� `�r߄ߖ�U���y��� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������	�� -��Tfx��� ����,> ��bt����� ��//(/:/��[/ /AC/�/�/�/�/  ??$?6?H?Z?l?~? �?O�?�?�?�?�?O  O2ODOVOhOzO�OK/ �Oo/�O�O�?
__._ @_R_d_v_�_�_�_�_ �_�_�?oo*o<oNo `oro�o�o�o�o�o�o �O�O�O5�O\n �������� �"�4��_X�j�|��� ����ď֏����� 0��o9]���I�� ��ҟ�����,�>� P�b�t���E�����ί ����(�:�L�^� p���A�S�e�w�ٿ��  ��$�6�H�Z�l�~� �Ϣϴ����ϗ����  �2�D�V�h�zߌߞ� �������ߥ���ɿ+� �R�d�v����� ��������*���N� `�r������������� ��&8��	�� }?������ "4FXj|;� ������// 0/B/T/f/x/�/I�/ m�/��/??,?>? P?b?t?�?�?�?�?�? �?�/OO(O:OLO^O pO�O�O�O�O�O�O�/ �O�/!_�/H_Z_l_~_ �_�_�_�_�_�_�_o  o2o�?Vohozo�o�o �o�o�o�o�o
. �OO_s5_7�� �����*�<�N� `�r���Co����̏ޏ ����&�8�J�\�n� ��?��cşן���� �"�4�F�X�j�|��� ����į֯������ 0�B�T�f�x������� ��ҿ��۟����)�� P�b�tφϘϪϼ��� ������(��L�^� p߂ߔߦ߸�������  ��$��-��Q�{� =Ϣ�����������  �2�D�V�h�z�9ߞ� ����������
. @Rdv5�G�Y�k� ����*<N `r������� �//&/8/J/\/n/ �/�/�/�/�/�/�� �?�F?X?j?|?�? �?�?�?�?�?�?OO �BOTOfOxO�O�O�O �O�O�O�O__,_�/ �/?q_3?�_�_�_�_ �_�_oo(o:oLo^o po/O�o�o�o�o�o�o  $6HZl~ =_�a_��_���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П����<�N� `�r���������̯ޯ ���&��J�\�n� ��������ȿڿ��� �"��C��g�)�+� �ϲ����������� 0�B�T�f�x�7��߮� ����������,�>� P�b�t�3ϕ�WϹ��� ������(�:�L�^� p���������������  $6HZl~ ���������� ��DVhz�� �����
//�� @/R/d/v/�/�/�/�/ �/�/�/??�!� E?o?1�?�?�?�?�? �?OO&O8OJO\OnO -/�O�O�O�O�O�O�O _"_4_F_X_j_)?;? M?_?�_�?�_�_oo 0oBoTofoxo�o�o�o �oO�o�o,> Pbt����� �_�_�_��_:�L�^� p���������ʏ܏�  ���o6�H�Z�l�~� ������Ɵ؟����  ����e�'����� ��¯ԯ���
��.� @�R�d�#�u������� п�����*�<�N� `�r�1���U���y��� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ���������	��� 0�B�T�f�x������� ����������> Pbt����� ����7��[ �������  //$/6/H/Z/l/+ �/�/�/�/�/�/�/?  ?2?D?V?h?'�?K �?�?�/�?�?
OO.O @OROdOvO�O�O�O�O }/�O�O__*_<_N_ `_r_�_�_�_�_y?�? �?�_o�?8oJo\ono �o�o�o�o�o�o�o�o �O4FXj|� ��������_ o�_9�c�%o������ ��ҏ�����,�>� P�b�!��������Ο �����(�:�L�^� �/�A�S���w�ܯ�  ��$�6�H�Z�l�~� ������s�ؿ����  �2�D�V�h�zόϞ� ���ρ������ɯ.� @�R�d�v߈ߚ߬߾� �������ſ*�<�N� `�r��������� ����������Y�� ���������������� "4FX�i� ������ 0BTf%��I�� m����//,/>/ P/b/t/�/�/�/�/� �/�/??(?:?L?^? p?�?�?�?�?w�?� �?�$O6OHOZOlO~O �O�O�O�O�O�O�O_ �/2_D_V_h_z_�_�_ �_�_�_�_�_
o�?+o �?OoOo�o�o�o�o �o�o�o*<N `_������ ���&�8�J�\�o }�?o����wڏ��� �"�4�F�X�j�|��� ����q֟����� 0�B�T�f�x������� m�����ۯ�Ǐ,�>� P�b�t���������ο ���ß(�:�L�^� pςϔϦϸ�������  ߿�	��-�W��~� �ߢߴ����������  �2�D�V��z��� ����������
��.� @�R��#�5�Gߩ�k� ������*<N `r���g��� �&8J\n ����u������ ��"/4/F/X/j/|/�/ �/�/�/�/�/�/�? 0?B?T?f?x?�?�?�? �?�?�?�?O��� MO/tO�O�O�O�O�O �O�O__(_:_L_? ]_�_�_�_�_�_�_�_  oo$o6oHoZoO{o =O�oaO�o�o�o�o  2DVhz�� ��o���
��.� @�R�d�v�������ko ͏�o�o�*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� ����C���|��� ����Ŀֿ����� 0�B�T��xϊϜϮ� ����������,�>� P��q�3��ߧ�k��� ������(�:�L�^� p����e�������  ��$�6�H�Z�l�~� ����a߫߅�������  2DVhz�� �������. @Rdv���� ���������!/K/ r/�/�/�/�/�/�/ �/??&?8?J?	n? �?�?�?�?�?�?�?�? O"O4OFO//)/;/ �O_/�O�O�O�O__ 0_B_T_f_x_�_�_[? �_�_�_�_oo,o>o Poboto�o�o�oiO{O �O�o�O(:L^ p������� �_�$�6�H�Z�l�~� ������Ə؏����o �o�oA�h�z����� ��ԟ���
��.� @��Q�v��������� Я�����*�<�N���o�1������$F�MR2_GRP �1a���� �C4  �B�[�	 [��߿�ܰE�� Fw@ 5W��S�ܰJ��NJk��I'PKHu���IP�sF!{���?�  W��S�ܰ9�<9��896C�'6<,5�{��A�  ��6��BHٳB�հ��޷�@�33�3�3S�۴��ܰ@UUT'�@��8���W�>u.�>*�߭<����=[��B=���=�|	<�K�<��q�=�mo����8�x	7H�<8�^6�?Hc7��x?��� �������"��F�X����_CFG b»T Q���|��X�NO º/
F0�� ��W��RM_CHKTYP  ��[�ʰ̰܂���ROM�_MsIN�[���9�u���X��SSBh��c�� ݶf�[�]����^��TP_DEF_O��[�ʳ��IR�COM���$G�ENOVRD_D�O.�d���THR�.� dd��_E�NB�� ��RA�VC��dO�Z�� ���Fs  G�!� GɃ�I��C�I(i J����+���%������ �QOUU��j¼������<6�i�C`�;]�[�C�հ��հȡ`��[�@ر����.��.R SMT��k_	ΰ�\��$HOST�Ch�1l¹[�̭d� 	�(�+��/Z��/W�e �/??'?9?G:�/j?�|?�?�?�/�?W0	anonymouy  �?�?	OO-O?N�/�/ �/�O�?�/Y?�O�O�O _K?(_:_L_^_p_�O �?�?�_�_�_�_ oGO YOkO}O_lo�O�o�o �o�o�o_�o 2 Dgo�_�_���� �o-o?o�S@��o d�v������o��Џ� ��)�*�qN�`�r� ���������� I�&�8�J�\�n����� ����ȯگ��3�E�"� 4�F�X�j���ß՟�� �ֿ�����0�B� �f�xϊϜϿ���� ������,�s����� ���߽�߿�������� �K�(�:�L�^�p�� ���ϸ������� �G� Y�k�}��l��ߐ��� ��������� 2 U�C��z�����//h!ENT 1m� P!V  7 ?.c &�J�n��� /�)/�M//q/4/ �/X/j/�/�/�/�/? �/7?�/?m?0?�?T? �?x?�?�?�?O�?3O �?WOO{O>O�ObO�O �O�O�O�O_�OA__ e_(_:_�_^_�_�_�_��ZQUICC0 �_�_�_?od1@oo.o�od2�olo~o�o�!ROUTER��o�o�o/!PC�JOG0!�192.168.�0.10	o�SCA�MPRT�\!bpu1yp��vRT�o���� !So�ftware O�perator Panel�mn���NAME !~�
!ROBO��v�S_CFG 1�l�	 ��Auto-st�arted'�FTP2��I�K2� �V�h�z������� ԟ����	���@�R� d�v���	������ �:���)�;�M�_�&� ��������˿�p�� �%�7�I�[��"�4� F�ڿ��������!� 3���W�i�{ߍߟ��� D���������/�v� �Ϛ�w�ߛ��Ͽ��� ������+�=�O�a� ��������������� 8�J�\�n�p�]�� �������� #5X�k}�� ��0/D1/ xU/g/y/�/RH/�/ �/�/�//?�/??Q? c?u?�?���/? �?:/O)O;OMO_O&? �O�O�O�O�O�?pO_ _%_7_I_[_�?�?�? t_�O�_O�_�_o!o 3o�OWoio{o�o�_�o Do�o�o�o����_ERR n���-=vPDUSIZW  �`^�P�Tt�>muWRD ?�΅�Q�  guest�f�������~�S�CDMNGRP �2o΅WpC��Q�`���fKL�� 	P01.0�5 8�Q   ��|��  };|��  z[� ���w����*���Ť�x����[ݏȏ�V�בPԠ���~���)����D�Yr���؊p"�P�l�P���Dx��d�x�*�����%�_GR�OU7�pLyN���	/�o���QUP���UTu� �T�YàL}?pTT�P_AUTH 1�qL{ <!i?Pendan�����o֢!KAR�EL:*������KC��ɯۯ���� ,��*�w�N�`����� ��㿺�̿޿+����X�CTRL r�L}O�uſa
�a?FFF9E3-ϝT�FRS:DEF�AULT��F�ANUC Web Server�� ��u�X���t@����1�C�U�g�;tWR_�CONFIG �s;� ��=qI�DL_CPU_P5C���aBȠP��w BH��MIN����q��GNR_IO�Fq{r�`Rx��NPT_SIM_DO���STAL_S�CRN� �.�I�NTPMODNT�OLQ����RTY�0����VIS\�E�NBQ�-���OL_NK 1tL{�p ������)�;�M���MASTE�%����SLAVE u�L|�RAMCAC�HEk�c�O^�O_�CFG������UO�C�����CMT_O�P���PzYCL�������_ASG s1v;��q
 O� r������� &8J\W�EWNUMzsPy
���IP����RTRY_CN��M�=�zs����Tu �������w���p/�p��P_�MEMBERS �2x;�l� $��X"��?�Q'W/i)���RCA_ACC �2y�  X��S�  ҿb6���"M����&6?��  H��/�(��%�(�$BUF00�1 2z�= �S�u0  u0�S��qP�Sf�:4g:4h:4i:4j�:4k:4l:4m:4n��<p�<q:4r:4s�:4t:4u:4v:4w�:4x:4y:4z:4{�:4|:4}L�:4��:4�:4�:4�:4��:4�:4�:4�RL��:4�:4�:4�:4��:4�:4�:4�:4��:4�:4�:4�:4��:4�:4�:4�:4��:4�:4�:4�:4�J:4�:4�:392$?�63P�.�A00�H1:1P1URY0URa0 URi0URq0URy0UR�0 UR�0�Z�0�Z�0UR�0 UR�0UR�0UR�0UR�0 UR�0UR�0UR�0UR�0 UR�0UR@UR	@j@ UR!@UR)@UR1@UR9@ URA@URI@URQ@URY@ ]ji@URq@URy@UR�@ UR�@UR�@UR�@UR�@ UR�@UR�@UR�@UR�@ UR�@UR�@UR�@UR�@ UR�@UR�@UR�@URP UR	PURPURP:193-_65WPA2WPI2WS NrY2gSNri2wSNry2 �SNr�2�x�2�x�2�S Nr�2�SNr�2�SNr�2 �SNr�2�SNr�2cNr 	B�B'cNr)B7cNr 9BGcNrIBWcNrYBh� iBwcNryB�cNr�B�c Nr�B�cNr�B�cNr�B �cNr�B�cNr�B�cNr �B�cNr�BsNr	Rs�NrR'v��2{�4(r�}ŋ���<����po�o��2�HIS!2�}� ܷ! �2024-07-	2� 1��П��� �ǹ!n��+�=�O�a� .�s�!������ί� ���(�:�L����� ��������ʿܿ� � �$�[�m�Z�l�~ϐ� �ϴ���������3�E� 2�D�V�h�zߌߞ߰� ������/��.�@� R�d�v������� �����*�<�N�`� r�������,P������@����#� o�c$ Oas������� ��'9K] o������� �/#/5/G/~�}/ �/�/�/�/�/�/�/? ?V/h/,?g?y?�?�? �?�?�?�?�?.?@?R? ?OQOcOuO�O�O�O�O �O�OO*O_)_;_M_ __q_�_�_�_�_��5p ������o$o6oHo� _oqo�o�o�o�o�O_ �o%7I[m ��o�o���� �!�3�E�W�i��� ����ÏՏ����� /�A�x����������� ��џ�����+�b� t�a�s���������ͯ ߯��:�L�9�K�]� o���������ɿۿ���I_CFG 2~��[ H
Cy�cle Time��Busy��Idl��mi�n�S�Up|��Read(ǟDowG�C� �W��Coun}t�	Num �"����� `����oPROG���U��P�)/so�ftpart/g�enlink?c�urrent=m�enupage,?1133,1�C��U�g�y�Tä�SDT�_ISOLC  ��Y� ���J�23_DSP_ENB  ��T���?INC ��� c���A   ?� � =���<#��
���:�o ��2�D� a/�l���OB��C��O��ֆ��G_GROUP �1���9d<�*�����t�?"���� `Q'�L� ^�p�/�����������\�~�G_IN_�AUTO����PO�SRE���KANJI_MASK0���DRELMONG ��[�� by�� ������f��%����� d-���KCL_L N�UM��G$KEYLOGGINGD��P�������LAN�GUAGE ��U��DE?FAULT ��Q�LG�����S��� ax�  �8T�H  � `'U0�� `; `�ލ�;��
*!(�UT1:\ J/ L/Y/k/}/�/�/�/ �/�/�/�/$>(�H?��VLN_DISP ���P�&�$�^4�OCTOL�0 aD�z����
�1GBO_OK ��d40V�11�0X,O !O3OEOWOiKyM�T��IgF	�5)�����O}���2_BUF�F 2��� � `2O�_�2��6_ M�R_d_�_�_�_�_�_ �_�_�_o3o*o<oNo�`o�o�o�o�o���ADCS ������ �L�O��+=Oa��dIO 2��kc +����� �������*� :�L�^�r��������� ʏ܏���$�6�J�~uuER_ITM��d������ǟٟ��� �!�3�E�W�i�{��� ����ïկ�����7Nx�SEVD��t�TYP����s���8���)RSTe�e�SCRN_FL +2��}���π�/�A�S�e�wϨ�T�P{��b��=NG�NAM��E��dU�PSf0GI��2�����_LOADދ�G %��%REQMENU����<MAXUALR�Mb2�@���
�K���_PR��2  h�3�AK�Ci0���qO=_'X�Ӭ�P 2]��; �*V	��-��
*����4 ��*��'�`�	xN�� z����������� 1�C�&�g�R���n��� ��������	��? *cFX���� ���;0 q\������ �/�/I/4/m/X/ �/�/�/�/�/�/�/�/ !??E?0?i?{?^?�? �?�?�?�?�?�?OO�AOSO6OwObO�OD�D�BGDEF ���գѢѤO�@_LDXDISA����ssMEMO_AP���E ?��
 �A�H$_6_H_Z_l_�~_�_�_K�FRQ_�CFG ���6�CA �G@��S�@<��d%�\o�_�P��Ґ�����*Z`/\b **:eb�DXojho�F �o�o�o�o�o�o ;�O��dZ�U�y|��z,(9�Mt� ��1��B�g�N��� r��������̏	����?�A�ISC 1���K` ��O���� �O���O֟����K�]��_MSTR ��3��SCD 1�]��l��{��� ��دïկ���2�� V�A�z�e�������Կ �������@�+�=� v�aϚυϾϩ����� ����<�'�`�K߄� oߨߓߥ�������� &��J�5�Z��k�� ������������� F�1�j�U���y����� ��������0T�?x�MK�Q��,��Q�$MLTA[RM�R�?g� ~s�@���@�METPU�@l���4�NDSP_ADCOL�@!oCMNT7 *�FNSW(FST�LIxi%� ��,����Q��*P�OSCF�bPgRPMV�ST5�1�,� 4�R#�
g!|qg%w/�'c/ �/�/�/�/�/�/?�/ ?G?)?;?}?_?q?�?��?�?�?�1*SIN�G_CHK  �{$MODA�S�e���#EDEV� 	�J	MC}:WLHSIZE�M�l �#ETASK �%�J%$123456789 �O��E!GTRIG 1�,� l�Eo#_`�y_S_�}�FYP�A��u9D"CEM_I�NF 1�?k�`)AT&FVg0E0X_�])�Q�E0V1&A3&�B1&D2&S0�&C1S0=�])�ATZ�_#o
dH@'oOo�QC_wohAo@�obo�o�o�o �_ &�_�_�_o�3o� �o���o��"�4� �X���ASe ֏���C�0��� f�!���q�����s�� ������͏>��b��� s���K���w���ٯ �ɟ۟L����#��� ��Y�ʿ����$� ߿H�/�l�~�1���U� g�y����ϯ� �2�i� V�	�z�5ߋ߰ߗ��߾PONITOR�G� ?kK   	?EXEC1o�U2�3�4�5�T�@�7�8�9o����(�� 4��@��L��X��@d��p��|��2��U2��2��2��2��U2��2��2��2��U2��3��3��3(��#AR_GRP_S�V 1��[ (0s��E�A_DsҔN~��ION_DB-@��1Ml  �bl #FH"4�l �FH��N BL6>FI-ud1}E����)PL_NA_ME !�E� ��!Defau�lt Perso�nality (�from FD)�b*RR2�� 1��L�XL�yp�X  d�� :L^p���� ��� //$/6/H/@Z/l/~/�/�/c2) �/�/�/??,?>?P?b?t?f<�/�?�?�? �?�?�?
OO.O@OROHdOc	�6�?�N
�O�OfP�O�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_�O�O2oDo Vohozo�o�o�o�o�o �o�o
.@o!o v������� ��*�<�N�`�r������ Fs  �GT�G�M�e���ÏՍfd�����(�6�������
��y�d����� ������ğ֟�� ���:���
�]�m�f��	`������į>��:�oAb	�����c A�  /���P����r� ������^�˿ݿȿ���%��R�� 1���	X ��, �� ��� a� @oD�  t�?�z��`�?f |�fA/���t�{	��;�	l���	 �xoJ����� �� �<�@����� ����K��K ��K=�*�J���J�?��J9���
�ԏC��@�t��@{S�\��(E�hє��.��I���ڌ���T�;f�ґ�$��3���´  �@���>�Թ�$�  >̿���ӧUf�g�x`���� ��
���Ǌ��� _�  {x @T�}����  �H ��l�ϊ�-�	'�� � ��I� �  �<��+�:�È��È�=�����x����N �[��n �@���f����f��k���,�av�  '���Yэ�@2��@�0@�Ш����C��Cb C���\C������G��@�� (�l�@X*�Bb $/�!��L��Dz�o�ߓ�~����( �� -���������!����D�  ��恀?��ffG�*<� !}�q��8���B�>��bp��(�(���P��	������>�?����x�����<
6b<���;܍�<����<���<�^���I/��A�{���fÌ�,�?fff�?_�?&� T�@��.�"�J<?�;\��"N\�3��� �!��(�|��/z��/j' ��[0??T???x?c? �?�?�?�?�?�?3��%F��?2O�?VO�/�wO�)IO�OEHG@� G@0��G�� G}ଙO�O�O_�	_B_-_f_Q_BL
��B��Aw_[_�_b� �_�[�_��mO3o�OZo��_~o�o�o�o���bs��PV( @|po 	lo-*cU�ߡ!A���r5eCP�xLo�}?�����#��3��W�s���6�Cv�q�CH3� j�t����q������|^(hA� ��ALffA]���?�$�?���;�°u�æ��)�	ff��?C�#�
����g\)�"�33C��
�����<��؎G�B����L�B��s�����	";�H�ۚG���!G��WI�YE���C��+�8�I۪�I�5�HgM�G�3E��R�C�j=x�
�p�I���G��f�IV=�E<YD�C<�ݟȟ�� ��7�"�[�F��j��� ����ٯį���!�� E�0�i�T�f�����ÿ ���ҿ����A�,� e�Pω�tϭϘ��ϼ� �����+��O�:�s� ^߃ߩߔ��߸����� � �9�$�6�o�Z�� ~������������ 5� �Y�D�}�h����� ����������
C:.(䁳��/"����<��xt��q3�8��<��q4Mgu����q�VwQ�
4p�+4�]$ $dR�v���u%PD"P��Q�_/�Z/=/(/a/L+R�g/n/�/�/�/�/�/  %��/�/+??O? :?s?/�_�?�?�?�;�?�?O�? OFO4O�rLO^O�O�O�O��O�O�J  2 {FsH�GT�V�M�uBO�|r�pp�C��S@�R_d_@v_�_�_�_�]�s\!�WɃooo�(o�z?���@@*�zh4�p�pk1u�p�~
 6o �o�o�o�o�o�o );M_q�ڊsa� ����D���$MR_CAB�LE 2��� ]��T��LaMa?�PMaLb�p�%Z��&P�C�p�!O4>�B]�%��~�v�l  ��&Py�v�wdN�{0�P��6�H�XT��6Pv� C$�Čj�(|����t ��&P��9C���=�о�Џ ��s9��T�,�>��� b�������Ɵ��Ο3� .��P�(�:���^�������������H�Z�l�*** �sOM ���y�����#%% 23�45678901�ɿ۵ ƿ���� ��� AQ� �!
��z�not s�ent ���W��TESTF�ECSALG� e�g;jAQd��ga%�
,���@���$�r�̹������� 9�UD1:\mai�ntenance�s.xmS�.�@��vj�DEFA�ULT�\�rGRP� 2���  p��Xwk  �%1�st mecha�nical chgeck��!���#������E��Z��(�:�L�^��"��c�ontrolleAr�Ԍ��߰��D������ ��$�s�M��L��""8b���v��B�����������/�C}�a�6����dv���s��C��ge��. b?attery�&��E	S(:L^�p�	|�duiz�awblet  D��"��R����/"/4/s��g�reas��'f�Br#-� |!�/�E�@�/�/�/�/�/s�
��oi,�g/y/�/��/t?�?�?�?�?s�H�
�XֈW��1<X�AO�E
c?8OJO\OnO�O�t��?O��'O�O_ _2_D_s��OverhaulE��L��R xX��Q�_���O�_�_�_�_oX�$�_0o����_o �_�o�o�o�o�o o�o?oQocoJ\ n���o�) ��"�4�F���|� �k��ď֏���� [�0�B���f������� ����ҟ!���E�W�,� {�P�b�t�����矼� ���A��(�:�L� ^�����ѯ㯸��ܿ � ��$�s�Hϗ��� ~�Ϳ�ϴ�������9� �]�o�Dߓ�h�zߌ� �߰�����#�5�G��� .�@�R�d�v��ߚ��� ���������*�y� ��`���O�������� ����?�&u�J�� n�����) ;_4FXj| ����%�/ /0/B/�f/���/ ��/�/�/�/?W/,? {/�/b?�/�?�?�?�? �??�?A?S?(Ow?LO ^OpO�O�O�?�OOO +O�O_$_6_H_Z_�O ~_�O�O�O�_�_�_�_po o�P�R	 T"o Ooaoso�_�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
���  ��Q?�w  @�a �o W�i�{��fC�����̟�h*�**  �Q�V��� �2�D��ph�z��������_ �S������կ7� I�[�����ɯ/���ǿ ٿ#���!�3�}��� ��{ύϟ��s����� ��C�U�g��S�e�w߀9ߛ߭߿�	�߉e��a�$MR_HI_ST 2��U��� 
 \jR$ �23456789C01*�2����)�9c_���R��a_�� �������=�O�a�� *�x�����r����� ��9��]o&� J�����# �G�k}4��d��SKCFMAPw  �U�)����`���ONREL  �����лEX_CFENB'
���!FNC$/$JOGOVLIM'qd�m �KEY'�p%y%_PANp(�"�"�RUN`,�p%�SFSP�DTYPD(%�S�IGN/$T1M�OTb/!�_C�E_GRP 1��U�"�:`��n? �c[?�?�؆?�?~?�? �?�?!O�?EO�?:O{O 2O�O�OhO�O�O�O_ �O/_�O(_e__�_�_ �_�_v_�_�_�_o����QZ_EDIT�4��#TCOM_�CFG 1���'%to�o�o 
Ua_/ARC_!"��O)�T_MN_MOD�E6�Lj_SP�L�o2&UAP_C�PL�o3$NOCH�ECK ?� � Rdv ����������*�<�N�`��NO_WAIT_L 7lJg50NT]a����UZ��_ERR&?12���ф��	� �-����R�d����`�O����|  ��
o��Z<� �� ?���ϟ�����ق_PARAMႳ���᠟R�g8�o��� = e ������گ�ȯ��"��4��X�j�F�g������A�ҿ�"ODR�DSP�c6/(OF�FSET_CAR8@`�o�DIS��wS_A�`ARK7�KiOPEN_FI�LE4�1�aKf�`O�PTION_IO��/�!��M_PRGw %�%$*��l��h�WOT��E7O����Z��G  �O�"�÷"�	 �W"��Z���RG_DS�BL  ���ˊ���RIENTkTO ZC����A �U�`IM�_D���O��V~�LCT ����Gbԛa�Zd��_�PEX�`7�*�RA-T�g d/%*���UP ���{��������������/$PAL�������_POS_CHU��7����2>3�L��XL�p��$�ÿU�g�y��� ������������	 -?Qcu����Y2C���" 4FXj|�� ���� //$/6/@H/Z/l/~/�Y�� �.��/�/ςP�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO�/ �/LO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_)O;O�_�_�_�_�_ �_�_o o2oDoVoho�zo�o�o�_����o�m ���~ BPw�m�m���~�jw#Ьw���� ��2�T��p��w���H��t	`���̏ޏ��:�o������ �2���A�   I��j�`������ ���џ���@���#�)�Or�1����� 8�>��, �\Ԡ�~� @D�  ��?���~�?� ���!�D������%G� � ;�	l��	 ��x�J젌����� ��<� ��� ���2�H(��H�3k7HSM5G��22G���GN�3%�R��oR�d��2�Cf��a��{���������/��3��-¸��4��>����𚿬���3�A�q�½{q�!ª��ֱ� "�(«�p=�2����� ��_{  @�Њ��_�  ��Њ��2��ς�	'� �� ��I� ��  �V���=�������˖ß���  �y��n @"��]�<߭�"��������N�Д߇  '�Ь�w�ӰC>��C��\C߰���Ϲ��ߤ!���@��4� (l~0�@X�B��B�I�;�)�j客z+���쿱����������( �� -��#�������!�]�9�|�  q�?�ffaH�Z��� ������"��8� ����>�|P$��}�(� ��P��������\�?���� x� ���<
6�b<߈;܍��<�ê<���<�^�*�gv�A)ۙ�脣��F��?fff?}�?&�� ��@�.���J<?�\��N\��)������� ����ޤy�N9 r]������ �/&/�J/5/n/��	g/�/c(G@� G@0i�G�� G}���/??<?�'?`?K?�?o?BL
i�B��A�?y?�?|� �?K�?ů�/QO�/xO��?�O�O�O�Om��bs��n�t @|�O '_�OK_6_H_�_lS��!A��RS�i�Cn_�_xj_0O�]?��o�oAo,où�Wi����ToC���`CH�Qo>Jd�`a�a@�Iܚ>(hA�� �ALffA�]��?�$�?����ź°u��æ�)�	ff���C�#�
ܢopg\)��3�3C�
������<��nG��B���L��B�s�����	0źH����G��!G���WIYE����C�+�½I�۪I�5�H�gMG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo�� �
��U�@�y�d��� ������я����� ?�*�c�N���r����� ���̟��)��9� _�J���n�����˯�� �گ�%��I�4�m� X���|���ǿ���ֿ ���3��W�B�Tύ� xϱϜ���������	� /��S�>�w�bߛ߆� �ߪ߼�������=��(�a�L�(q���)����Z�������a3�8�������a4Mgux�����a�VwQ��(�4p�+4�]B�B���p�����������UPbP���Q O%x�1[FjR�������  C���I 4mX�8
O������.//>/d/R/�Rj/|/�/�/�/�/�/:  2� Fs�gGT]�&6�M�eBmpX�R�P�aC��3@�_ p?�?�?�?�?�?�=�S�OO)O;OMO�c�?���@@�jJ��`�`�1�`�^
 TO�O�O �O�O�O_#_5_G_Y_�k_}_�_�_�j�A �����D��$�PARAM_ME�NU ?B���  �DEFPULS�E�[	WAIT�TMOUTkR�CVo SH�ELL_WRK.�$CUR_STY�L`DlOPT�Z1ZoPTBooibC�?oR_DECSN `���l�o�o�o &OJ\n������QSSREL_ID  >��
1��uUSE_P�ROG %�Z%8�@��sCCR` ��
1�SS�_HOST7 !�Z!X����M�T _���x�������L�_TIME�b �h��PGDE�BUG�p�[�sGI�NP_FLMSK��E�T� V�G�PG�Ar� 5��?��CyHS�D�TYPE�\�0��
�3�.� @�R�{�v�����ï�� Я����*�S�N� `�r����������޿ ��+�&�8�J�s�n���ϒϻ�G�WORD� ?	�[
 	�PR2��MA9I�`�SU�a��cTEԀ���	Sd�COL��C߸��L� C�~��h�d*�TRACE�CTL 1�B�]�Q ��0�'�߫Ӂ�DT Q�B��М�D 7� ������ ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OE�� .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� "Op���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| �d������ 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o��o�o�c�$PGT�RACELEN � �a  ����`��f_�UP ���e�q'pq   p��a_CFG ��u	s�a p��LtLtfqwpqz�  �qu4rDEFSPD �?|��ap��`H_�CONFIG ��us �`j�`d�t��b �a��qP�t�q��`���`IN7pTRL ��?}_q8�u�P�E�u��w��qLt�qqv�`LID�8s�?}	v�LLB� 1��y 5��B�pB4Ńqv �އ؏	�s� <<0p  ?��'���A� o�U�w�������۟���ӟ��#�	�+�Y�v� 񂍯����ï
���������/�u�GRP �1ƪ��a@俼j��hs�aA��
D�� D�@� Cŀ @�٭^�t�q�����q�p���.� ���FȾ´���ʻB� )�	���?�)�c��a�>��>�,���Ϻ��ζ� =49X=H�9��
��� �@�+�d�O���s߬��o߼�����  Dz���`
��8���H� n�Y��}������� ������4��X�C�|����)��
V7.10beta1Xv A�������!�����?!G��>\=y��#��{33A!�ߚ@��͵��8�wA��@� A�s�@Ls���� ��"4FXLsAp,ry��q��� ��q�ar�T�n�t�����	t�KNO?W_M  |uGv�z�SV ��z�rs&����>�/�/G/�a��y�M�M���{ ���	~^u (l+/��/',_t@%X�����@���%��"4�.0pz�MR
M��|-TU�y�c?�u;eOADBANgFWD~x�STM��1 1�y�4e��8��̾�?�?�? (OO-O?OqOcOuO�O �O�O�O�O�O&___ \_;_M_�_q_�_�_�7�2�<�!�?�`�<�_�_N�3�_�_
oo��749oKo]ooo�75 �o�o�o�o�76�o�o�772DVh��78�����7M�A�0��swwO�VLD  �{��/a�2PARNUM  �;]�o��3�SCH*� 8�
�����ω�3�UPD���[�ܵ+�wu_CM�P_r -��0�'��5C�ER_CHKQ����1�"e�N��`�RS>0�?G�_M�O�?_��#u_R�ES_G�0��{
 Ϳ@�3�d�W���{� �������կ���*� ����P��O� �8`l�������`�� ʿϿ��`�	��� 1p)�H�M���phχπ����p�������V� 1��5�1�!@�`y�ŒTHR_�INR>0/�Z"�5d�:�MASSG� Z�[�MNF�y�MON�_QUEUE ���5�6Ӑ~#tN�H�U��N�ֲ���E�ND�����EXE�����BE������OPTIO�������PROGRAM %��%��߰�~��TASK_I,��>�OCFG ��ߞ�����DATA�u#�����Ӑ2 �%B�T�f�x���5��� ����������,>�P�INFOu#� �������� �'9K]o ��������h/lx� � ;�l��ȀK_������S&ENB-�b-&q҂&2�/�(G��2��b+ X,		ޖ�=����/��@��P4$�0��9�9)�N'_EDIT� ���W?i?��W�ERFL�-ӱ3RGADJ �F:/A�  �5?Ӑ�5�Nј6��]!֐���?�  B�z�WӐ<1Ӑ�%��%O�8;��50!2ج�7�	H��l0��,�BP�0㎹@�0�M*�@/�B **:�B�O�F$�O2��D��A�ЎO��@O	_,X��%���H�q��O$_r_0_�_���Q@WA��>]�_ �_�_o�_o�_�_
o �o.o�ojodovo�o�o �o�o�o�o\XB <N�r���� 4��0���&���J� ������������� ���x�"�t�^�X�j� 䟎���ʟğ֟P��� L�6�0�B���f����� ����(�ү$���� ��>���z�t��� Ϫ� �����l��h�R�L�^�DX	���ώ0��< ���t$ :�L���o�
ߓߥ��7PR�EF ��:�0��0
�5IORIT�YX�M6��1MPD�SPV�:
B �UT���C�6ODUCT���F:��NFOG[@_TG�0��J:�?�HIBIT_D�O�8��TOENT� 1�F; (!AF_INE*������!tcp|���!ud��~8�!icm'���N?�XY�3�F<��1)� �A�����0��������� ��' ]D�h�������*>��3��9
BOTfN�3>���2�B�G!/�LC��4�;LFJ�AB,  � ��F!//%/7/�5�F�Z�w/�/�/�/��3&ENHAN�CE �2FBA�H+d�?�%;��������Ӓ1�1POR_T_NUM+��0����1_CAR�TRE�@��q�S�KSTA*��SL�GS�������C�Unothing?�?OO����0TEMP ��N�"O�E�0_a_?seiban|߅O xߕO�O�O�O�O_�O '__K_6_H_�_l_�_ �_�_�_�_�_�_#oo Go2okoVo�ozo�o�o �o�o�o�o1U @e�v���� �����Q�<�u�>.IVERSI	�L���� dis�able�.GSA�VE �N�	�2670H771|�h��!�/��9�:� 	^�4�ϐ�	���e��͟ߟ�����9�D�C-Å]_y� 1������ő����Ǻ�/URGE� B��r�WFϠ��-��9��W����l:WRU�P_DELAY ��=n�WR_HOT %��7��/�p��R_NORM�ALO�V�_�����S�EMI��������Q/SKIPo��97��xf�=�b�a�sυ�H� �ʹ��ø�������� &��J�\�n�4�Fߤ� �������߲���� � F�X�j�0��|���� �������0�B�T� �x�f���������ãRBTIF�5���CVTMOU�7v�5���DCRo�}�� �T��+댹^�Cj�P>�4J^�9L��&H�  �j=W�ſE���V�����<
6b<�߈;܍�>u�.�>*��<ȃ�ǪP0�� �2DVhz��������,GRD�IO_TYPE c v��/ED� �T_CFG �l�-�BH]�EP)v�2��+ ��B�u �/�*��/� ?�/%?=�/V?�}? �Ϟ?���?�?�?�?�? O
O@O*Gl?qO��8O �O�O�O�O�O�O�O�O _<_^Oc_�O�__�_ �_�_�_�_o�_&oH_ Mol_o�oo�o�o�o �o�o�o�o"DoIho *j����� ��.3�E��f� � ��x��������ҏ� *�/�N��b�P���t� ����Ο��ޟ�:�+����R'INT 2��R��!�1G;� �i�{��"���8f�0 ��ӫ���� ��M�;�q�W����� ��˿���տ�%�� I�7�m��eϣϑ��� ��������!��E�3� i�{�aߟߍ��߱����������A���EFPOS1 1�!)?  x��� n#����������� ��/��S���w���� 6�����l������� =O����6��� V�z� 9� ]����Rd ���#/�G/�k/ /h/�/</�/`/�/�/ ??�/�/?g?R?�? &?�?J?�?n?�?	O�? -O�?QO�?uO�O"O4O nO�O�O�O�O_�O;_ �O8_q__�_0_�_T_ �_�_�_�_�_7o"o[o �_oo�o>o�o�oto �o�o!�oEW�o >���^��� ��A��e� ���$� ����Z�l�����+� ƏO��s��p���D� ͟h�񟌟�'�ԟ �o�Z���.���R�ۯ v�د���5�ЯY��� }���*�<�v�׿¿�� ��Ϻ�C�޿@�y��e�2 1�q��-� g�����	��-���Q� ��N߇�"߫�F���j� �ߎߠ߲���M�8�q� ��0��T����� ���7���[����� T�������t�����! ��W��{�: �^p��A �e �$��Z �~/�+/��� $/�/p/�/D/�/h/�/ �/�/'?�/K?�/o?
? �?.?@?R?�?�?�?O �?5O�?YO�?VO�O*O �ONO�OrO�O�O�O�O �OU_@_y__�_8_�_ \_�_�_�_o�_?o�_ co�_o"o\o�o�o�o |o�o)�o&_�o ��B�fx� �%��I��m���� ,���Ǐb�돆���� 3�Ώ���,���x��� L�՟p�������/�ʟ�S��w�����ϓ�3 1��H�Z���� ��6�<�Z���~��{� ��O�ؿs����� ϻ� Ϳ߿�z�eϞ�9��� ]��ρ���߷�@��� d��ψ�#�5�G߁��� ����*���N���K� ����C���g���� �����J�5�n�	��� -���Q��������� 4��X��Q� ��q��� T�x�7�[ m�//>/�b/ ��/!/�/�/W/�/{/ ?�/(?�/�/�/!?�? m?�?A?�?e?�?�?�? $O�?HO�?lOO�O+O =OOO�O�O�O_�O2_ �OV_�OS_�_'_�_K_ �_o_�_�_�_�_�_Ro =ovoo�o5o�oYo�o �o�o�o<�o`�o Y���y� �&��#�\�����ए?�ȏ����4 1�˯u�����?�*�c� i���"���F����|� ���)�ğM����� F�����˯f�﯊�� ���I��m����,� ��P�b�t������3� οW��{��xϱ�L� ��p��ϔ�߸����� �w�bߛ�6߿�Z��� ~�����=���a��� �� �2�D�~������ ��'���K���H���� ��@���d��������� ��G2k�*� N����1� U�N��� n��/�/Q/� u//�/4/�/X/j/|/ �/??;?�/_?�/�? ?�?�?T?�?x?O�? %O�?�?�?OOjO�O >O�ObO�O�O�O!_�O E_�Oi__�_(_:_L_ �_�_�_o�_/o�_So �_Po�o$o�oHo�olox�oۏ�5 1��� �o�o�olW��o� O�s���2�� V��z��'�9�s�ԏ ���������@�ۏ=� v����5���Y��}� ����۟<�'�`����� ���C���ޯy���� &���J����	�C��� ��ȿc�쿇�ϫ�� F��j�ώ�)ϲ�M� _�qϫ����0���T� ��x��u߮�I���m� �ߑ��������t� _��3��W���{��� ���:���^����� /�A�{����� ��$ ��H��E~�= �a�����D /h�'�K� ��
/�./�R/� �/K/�/�/�/k/�/ �/?�/?N?�/r?? �?1?�?U?g?y?�?O �?8O�?\O�?�OO}O �OQO�OuO�O�O"_t6 1�%�O�O _�_�_�_�O�_|_o �_o;o�__o�_�oo �oBoTofo�o�o% �oI�omj�> �b������ �i�T���(���L�Տ p�ҏ���/�ʏS�� w��$�6�p�џ���� �����=�؟:�s�� ��2���V�߯z����� د9�$�]�������� @���ۿv�����#Ͼ� G�����@ϡό��� `��τ�ߨ�
�C��� g�ߋ�&߯�J�\�n� ��	���-���Q���u� �r��F���j���� ��������q�\��� 0���T���x����� 7��[��,> x����!�E �B{�:�^ �����A/,/e/  /�/$/�/H/�/�/~/�?�/+?�/O?5_GT7 1�R_�/?H?�? �?�?�/O�?2O�?/O hOO�O'O�OKO�OoO �O�O�O.__R_�Ov_ _�_5_�_�_k_�_�_ o�_<o�_�_�_5o�o �o�oUo�oyo�o�o 8�o\�o��? Qc���"��F� �j��g���;�ď_� 菃������ˏ�f� Q���%���I�ҟm�ϟ ���,�ǟP��t�� !�3�m�ί��򯍯� ��:�կ7�p����/� ��S�ܿw�����տ6� !�Z���~�Ϣ�=ϟ� ��s��ϗ� ߻�D��� ���=ߞ߉���]��� ��
���@���d��� ��#��G�Y�k��� ��*���N���r��o� ��C���g������� ����nY�-� Q�u��4��X�|b?t48 1�?);u��/ ;/�_/�\/�/0/ �/T/�/x/?�/�/�/ �/[?F???�?>?�? b?�?�?�?!O�?EO�? iOOO(ObO�O�O�O �O_�O/_�O,_e_ _ �_$_�_H_�_l_~_�_ �_+ooOo�_soo�o 2o�o�oho�o�o�o 9�o�o�o2�~� R�v���5�� Y��}����<�N�`� ��������C�ޏg� �d���8���\�埀� 	�����ȟ�c�N��� "���F�ϯj�̯��� )�įM��q���0� j�˿��ￊ�Ϯ�7� ҿ4�m�ϑ�,ϵ�P� ��tφϘ���3��W� ��{�ߟ�:ߜ���p� �ߔ���A����� � :����Z���~�� ���=���a���� ������MASK +1�������~��XNO  ����� MOTE  ��R_CFG ��Y����PL_RANGUP����OWER ���� �A���*SYSTEM*�P�V9.3044� �1/9/2020 A � ����RESTA�RT_T   �, $FLAG�� $DSB_S�IGNAL� $~UP_CND4����RS23�2r � �$COMMENT� $DEV�ICEUSE4P�EEC$PARI�TY4OPBIT�S4FLOWCO�NTRO3TIMgEOUe6CU�=M4AUXT��5�INTERFAC�sTATU���KCH� t $OL�D_yC_SW �'FREEFR�OMSIZ �A�RGET_DIR� 	$UPD�T_MAP"� T�SK_ENB"E�XP:*#!jFA�UL EV!�R�V_DATA�_  $n E��   	$VAL�U�! 	j&GR�P_   �{!A  2 ��SCR	�� �$ITP_��" $NUMΞ OUP� �#TO�T_AX��#DS}P�&JOGLI�FINE_PCdn�OND�%$�UM�K5 _MIiR1!4PP TN?8�APL"G0_EX�b0<$�!� 814�!P=Gw6BRKH�;&{NC� IS �  �2TYP� �2�"�P+ Ds�#;0BS�OC�&R N�5DU�MMY164�"S�V_CODE_O�P�SFSPD_�OVRD�2^L�DB3ORGTP; LEFF�0<G� �OV5SFTJRUNWC!SFpF5%3oUFRA�JTO��LCHDLY7R�ECOVD'� WaS* �0�E0RO���10_p@  � @��S NVE�RT"OFS�@C� "FWD8A�D4A��1ENABZ6�0T�R3$1_`1FD}O[6MB_CM�!zFPB� BL_M��(!2hRnQ2xCV�"�' } �#PBGiW|8A�Mz3\P��U�B�__�M�P�M� �1�AT�$CA� �PD�2��PHBK+!:&aI�O�4 eIDX+bPPAj?a$iOd�7e�U7a�CDVC_DBG"�a;!&�`��B5�e1�j�S�e3��f�@ATIO� ���AU�c� �S�AB
0Y.#0�D���X!� _�:&S�UBCPU%0S�IN_RS�T, 1�N|�S�T!�1$HW_C1�"]q.`�v��Q$AT! � �_$UNIT�4�p>�pATTRI= �r�0CYCL3NE�CA�bL3FLTR_2_FI9a7�c�,!LP;CHK�_�SCT>3F_ƥwF_�|8��zFS8+�R�rCHAGp�py��R�x�RSD�@`'�1E#&7`_T�X�PRO�`@S�EMOPER_0�3Tf��]p� f��P�DI�AG;%RAILAiC�c4rM� LO�04�A�65�"PS�"�2� -`�e�SPR�`S&.  �W�Ctaf�	�CFUNC�2~�RINS_T.!`(�w��� S_� ��0�P�� 	d��W�ARL0bCBLCUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!��8�3�TID�S��!�� $CE_RIYA !5AFDpPC�~��@��T2 �C�9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@HRgDYOL1	PRG8��H��>1(�ҥMUGLSE =#Sw3��$JJJ6BKGFK�FAN_ALML�V3R�WRNY�HGARD�0+&_P "B��2Q���!�5_�@�:&AU�Rk��TO_SBRvb��� �ƺ�pvc�޳MPINF�@�q�)���'REG'd~0V) 0R<�C�1DAL_ \2sFL�u�2$MԐ (�#S��P� `�gśCMt`NF�qsO�NIP�qEIPPs 9a$Y���!��"�!7� �o3EGP��#�@��AR� �c�52p�����|5AXE�'wROB�*RED�&�WR�@�1_=��3S�Y�0ѥ0_�Si�WcRI�@�ƅpST@�#��0*@� �q	���3��� B� �A��3�]D�POTO�� �@ARY�#��!��d̒!1FI�0�$�LINK��GTH��B T_���Ar��6�"/�XYZ+":9�7G�OFF�@�).�"���B� l�����A3$ ��FI@�p���4�4l��$_Jd�"(B�,a������8�"q�����2�Ck6DUR��]94�TURT�XZ��N����Xx��P��FL/�@s��l�P���30�"Q 1J� K
0M:$�53]q�7�SuD�Sw#ORQ�Ɇ�!�����Q7��0O[�ND�=#�!#�1'OVE8��M� ��R��R��Q!P0.!P! OAN}q	� R����990� �br J9V����v�!SER1��	8�E�@Hn D�A��p�����Ă���v�AX �C�"��`�q�s� ��0~3�~F��~e�~�~E�~1 ��~Ҡ{Ҡ�Ҡ� Ҡ�Ҡ�Ҡ�Ҡ��Ҡ�Ҡ�!)DEBU}s$x�����!R*�AB�a8Ar2V`|r 
�" �c���%�Q7�7�1 73�7F�7e�7�7E�������L�AB����yp�cG�RO�p��}��PB_ҁ ��̓��ð�6��1���5���6AND ��8p�a3���-G �Q����AH�PH�p�2�NTd��Cs@VE�L؁�}A��F�S�ERVEs@�� i$����A!�!�@POR}�KP�иA����@���	  �$�BTRQ�
��CH��@
�G��2	��Eb��_  qlb��Q�ERR��RI�P�@�FQTO	Q�� L�}��YV
ĀG�E%�\���B�RE�  ,h�A�EP
�RA�Q? 2 d�R7cs�T�@ ���$F ׂ��m  ��COC��P � 8[COUNT����@�PFZN_C;FG�A 4�p%��rT\zs�a�#`pJpx c%d�� �� MGp+����`�OGp��eFAq����cX�8еk�ioQ��'ѴD�p8�Pz���HEL�A�-b 5���B_BAS\RSSR$�`�2�S�ѤL�!p1�W!p2Dz3�Dz4Dz5Dz6Dz7rDz8�WqROO��P�1�NL�� �AqB�C
�"pACK�&KIN�PT+�W�U��8	�k��y_PU8�~�|�OU�CP��%�s��Vl���YTPFWD_KARKQ-�:PRE�D�P����QUE$�Ā9 )���~���IU��#s/��8�@�/�SEM1ǆt1�A�aSTY�t3SO����DI�q��pQc��X��_TM9ßMANRQ �/�E�ND��$KEY?SWITCH2�G�����HE)�BEA�TMz�PE��LEPJR���0x�UF�F���G�S�DO_HOeM��Oz��pEF�PR��SbJі��uC⒐O��7P�QOV_�M��}�c�IOCM����1�BsHK��� D,�&�a`U�2R��M��a�r +�FwORC*�WAR��hbsOM�� � @�$�㰰U��P��1��g���3��4��1�B�POW�Lz�<�R%�UNLO�0T��ED��  ��SNP��S.b; 0N�ADDa`z��$SIZ*�$�VA�0�UMULTKIP�r���Az� � $���ƒ���SQc�1C<FPv�FRIFr�PaSw���ʔf�NF#�ODBUx�R@w���0���F��:�IAh��Ƙ�������S"p��� �  �cRTE����SGL.�T�x�&C`Gõ3a�/�OSTMT��`�P����BW9 0�SHO�Wh�qBANt�TPo���E�������@V_Gsb �$PC�0�PokFBv�P��SP��1A�p���PVD��rb�� �+QA002D.ҝ�6ק�6�P��6׻�6�54�64�U74�84�94�A4�B4و�6ׇ17�}�6�F4� ��@�����Z٨���t�1��1��1���1��1��1��1���1��1��1��2�3�2@�2M�2Z�2�g�2t�2��2��2���2��2��2��2���2��2��2��3P3����M�3Z�3g�U3t�3��3��3��U3��3��3��3��U3��3��3��43�U4@�4M�4Z�4g�U4t�4��4��4��U4��4��4��4��U4��4��4��53�U5@�5M�5Z�5g�U5t�5��5��5��U5��5��5��5��U5��5��5��63�U6@�6M�6Z�6g�U6t�6��6��6��U6��6��6��6��U6��6��6��73�U7@�7M�7Z�7g�U7t�7��7��7��U7��7��7��7�ٕ7��7��7��#bV�Pv�U�B ��@�09r
Ѱ��A/ x �0R���+  �BM�@RP�`�4Q_�PR�@[U�A�R��DSMC��E�2F_U��=A�QY�SL�P�@ �  �ֲ>g�����x��iD��VALU>e��pL�A�HFZAID�_L���EHI�JI~h�$FILE_ ���D�d$ǓUFSA��Q h�0!PE_BLCKz�.RI�>7XD_CPUGY!� GY�Ic�O
TVA����R  � �PW`�p���QLAn�S�Q�S�Q�TRUN_FLG�U �T�Q�TJ��U�Q�T�Q��UH��T`�ThaT�2L�_LIz� w �pG_O}T�P_EDIU�-b�`7c ?bة�p�BQh�����TBC=2 �! �%�>�0�P��a�7aFTτ�d.݃TDC�PA�N`��`M�0�f�a�gTHD��U��d�3�gR�q<�9�ERVEЃt�݃t	��a�p�` "X -$EqLENЃRt݃Ep�pcRAv��Y@W_A�tS1Eq�D2�wMO$?Q�S���pI�.B`�A�y�4Ep�{DE�u���LACE �CCqC�.B��_MA�p�v��w�TCV�:��wT,�;�Z�P�Ҡ�s�~��s�J�A�M����J���u)ā�uQq2ѐ����݁�s�JK��V�K������	���J�����JJ�JJ�AAL�<��<��6��:�5�cm�N1�a�m�,��DL�p_x\�Ű,bBCCF
��# `�0GROUP�@J�Բ��N�`C^�~ȐREQUIRr�ÀEBUu�Aq��$T�p2"��Bp�8�a	��d$ \?@qhoAPPR��CLB�
$H`N;�CLOD}`K�S�e`��u
�a.I�% �3�M�`�8l��_MG񱥠�C �"P����&���B{RK��NOLD����RTMO6a�ޭ��J6`�P>��p���p��pZ��pc��p6�+�7+�<�	 |@r�d&� ��lr��������PATH��������qx��䋠�%0A��SCA�ub��<���INDrU�C�p�q�C�UM�Y�pP����A� q/ʤ�/�E�/�PA�YLOA�J2L��0R_AN�ap�L��Pz�v�jɆ���R_?F2LSHRt��LO{�R�������ACRL_�q������b�d�H�@B$yH��"�FLEX>�u�aJ�f' P(� �o�o+�p>�Du( :Qcv�p ����fe��po��|F1���-������]�E��*� <�N�`�r�����4�Q� ������A�c���ɏۏ$���T��2�X:A;� �������� )�;�?�H�6�Z�c�u�p����>Ѭ�) ��``��˟ݟ�`�0ATF�𑢀EL��(a���J�(��JE۠C3TR��A�TN�1��HAND_VB�B>ѯ@�* $���F2���d�CS�W>�����+� $$M�����0ˡ��ڡ������A@�@g����A)��A���@˪A٫A� ��T`P˪D٫D�PȰG�P�)STͧ�!ک�!N�DY�P9��� �#%��Fp���Ѫ���@i����������P3� <�E�N�W�`�i�r����e, ��ԓ� �n�5m��1ASYIMص.@�ض+A������_`��	�� �D�&�8�J�\�n�Ju�&��ʧC�I��S�_VIo�Hm��@V_UNVb�@
S+��J�"RP5"R��&T ��3TWV�͢���&��ߪU��/�7�=r�`3HR`ta-��QLQ�1�DI��O�T8���P��. ; *"IAA*���$aG�2C�2cJ��`y�I��P �/ � �MEB�� Mb�R4AT�PPT�@� ��ua���AP�l@zh�a�iT�@��� $DUM�MY1E�$PS�_D�RFॐ$��f3�FLA��Y�P���b}c$GLB_T��Uuu`1�p=Ѓ�EQa0 X(����ST����S�BR�PM21_V���T$SV_ERb��O_@KscsCLp�KrA��O'b�PGLv�@EW��1 4���a$Y|Z|W�s怯��AN`¼��qU�u2 ��N��p�@$GIU}$�q �p�s�p���3 L���v^B}�$F^BE�vNEA�R��NK�F8���T�ANCK����JO�G��� 4��?$JOINT����t�qMSET��5�  �wE�H�� S������ ��6�k  MU��?���LOCK_FO�����PBGLVHG�L�TEST_X9M>���EMPt���q�r̀$U�Ќ�r��22���s,�3����Ҁ,�1MqCE����sM� $KAR���M�STPDRA8�pj�a�VEC��{��e�IU,�41�HE�ԀTOOL㠓Vv�RE��IS3��r��6N�A�ACH����5��O�}c�d3ڲ��pSI.� � @$RAIL_�BOXE��ppR�OBO��?�pqHOWWAR*���`�ROLM�bB����S��
�5���O_�F� !ppHTML5�Q����С2�pڑ��7m��R��O��8���v��z���uOU��9 tpp(�14A��̀��PO֡%PIP��N��
�ڑ�S�,�����CORD�EDҀް̠5�XTT��q)bP� O4` : D pOBP!"Ҁ{�j��cppj�^@$SYSj��ADR#�Pu`TC}H� ; ,��SEN�RZ�Aف_�t�״��J`PVW�VAPa< � �p��r�UPREV�_RT]1$ED�IT�VSHWRB�7v;���q�@�D_`#R�+$HEADoA�Pl�A�$�KE�q�`CPwSPD��JMP��=L�U �TR��d�=r�O�϶I�S#CiNE��$_OTICK�AMX���Q��HN-q>� @t������_GqP��[�STYѲ�LOq�s��Ҩ��?�
�Gݵ%$����t=7pS !�$Q��da�e!`�fP�0�SQUd� ��b��ATERCy`�2�{TS�@ �p�Cp����d�%Oz`mcO�IZ�d�q�e�aPRM��a8�����PUQH�_DO�=�ְXS��K�VA�XIg�f�1�UR � ��$#�Е��� Y_����ET��Pۂ@���5�o��6g�A�!V�1�d9�2;�]�TSR|Al�о���#�� 5��#��#�)#�) i�>'i�N'i�^&{��� �){����2��C�����C��WOiO{O�DtS�SCp B h�ppDS(�k��`SPL`�ATL �I����¼bADDRE�S��B'�SHIF���"�_2CH#r��I&p��TU&p�I� C��CU�STO���QV��I�bDȲ,��0
��
z�U�R`E 	\�����f�7��tC�#	���F��ir�t�TXSCRE�El�F�P��TICNA�s�p��t��8���0G T��fp ,⧱eqBp&uᦲu�$#�RRO'0R����}�!����UE��H# ��0���`S�q��'RSM�k�UV����V~!�PS_�s�&C �!�)�'C��Cǂz"�� 2G�UE©4Ibvr�&8�GMTjPLDQ��Rp�^��BBL_�W�`NR`J �f�>2O�qJ2LE�U3"��T4RIGH^3BRyDxt�CKGR�`�5TW��7�1WIDTH�H������a��� �UIu�EY��QaK d�p��A��J�
�4�BACK�H��b�5|qX`FO�D�GLABS�?(�X`I�˂$UR�(�9@���0^`H4! OL 8�QR�_k��\B_`R�p͂���H�a^�IAO�R`M�I�w0Uj0�CRۂ�M�LUM�C��� E#RV��0P<��45NV`��GE=B#����]�t�LP�E��E��Z)Wj'Xz'XTԐ&Y5$[6$[7$[8	R���3�<���fjԑŁS��M�1�USR�tO <ļ�^`U�r�rFO\
�rPRI��m�����PTRIP��m�UNDO��P�p��`m�4�l�p�@$���� QWB\�P7�G s�Tf��H�RbOS�agfR ��:">c��.qR��s �~�b*��A$�UQ.q�S�o�o�#R)�>cOSFF���pT� �c=Op 1R�tZ/tS�GU��P.q๢JsETw�1SUB�*� f�E_EXeE��V��>cWO>� U�`^g��WQA'��P�q!@� �V_DB�s�p�BSRT�`
�V�Q�r���OR��uRAUD��tT�ͷ�q_�β�W |%�͸OW�NA`޴$SRC�E � ��D��\��M�PFIA�p��ESPD������C���G�ƒ)�5��!X `��`�r޴��COMP�a$��C`_w�`�����rCT�3 �q���qƒ��@�� Y"SHAD�OW�ઓ@�_UN�SCA��@��4M�D�GDߑ��EGAC��,Me�G�Z (0NO�@�D<�kPE�B��VW�� �G���![ � ���VEE#�aڒANG�$��c薴cڒLIM_X�c��c � ����#��`� ���bVF� �s�VSCCjв�\ՒC{ЃRAlצ���RpNKFA��%�E���Z`G� ^0[��C`DEĒ��� STEQ1���@�ꁻ@ I��`+0����`����P_A6�r���K�|���!]� 1�������\��сCP9C�@]�DRIܐ\�B͑V#Ѐ���D�T?MY_UBY�T��@�c��F!���Y�브����P_V�y��L�N�BMQ1$��DEY��EX�e���MU��X�M� U1S�!���P_R��b��P� ߖG��PACIr�ʐf�ᔟ��c���c���#�EqB��a�.2B����^ ܀GΐP���)�D�R~``�_�0�@3!��1zr	�e�R�S�W��p�00��S�6�OD�Q�1A� X�#�E��UE��00�HK
J�`�@p���U� �EAN�ٖp�pxXՆ`C�MRCV�!Wa ��@O��M�p�C�	��s����REF*7
�������� /��P��@���@��b��֗�_Y��ژ��ۣ� �Q$3������AC��$b ����%����Q��$GROU@� �c�����ʠ]��I2^0��U` 0�_�I,�o � U�Lա`��C&�rAaB�?�NT������@���A���Q��K�L�����õ��A���Q��T� a$c t�`MD��p8�HU���S]A�CMPE F(  _�Rr�p�@����XS	qVG�F/�b#d, &��@M�P^0۰UF_`C !���z �ROh0�"+���@���0C�UcREB���RI��
IN�p�����`d��d��ca�INE�H�y��0V�a-����3�W������0�C��i�LO�}��z�@0�!�QNSI ��݁���c$&�c$&.��X_PE-YW+Z�_M�ڒW�I��$�" �+R�'rRS�Lre �/�M�
`�RE�C7�G d�۰�̵ҭ�q���� u��Ȑ�������S_P�VnP *�I�A�vf �~pHD5R�p�pJO�P���$Z_UPz��a_LOW�5�1J�dA��LINubEP?�tc_i�1�1���@�G1@��V�x�g 5X�PA�THP X�CACH$�]E��yI�AT��{�C)�ID3FA�ETD�H��$HOD�pO�b@�{�d6��F�����p�PAGE�䁀VP�°�(RO_SIZ��2TZ3�`-X�0U�q�MPRZ���IMG���A9D�Y�MRE��R�7WGP��8�p��A�SYNBUF�V�RTD�U�T7Q�LE_2D-��U��`%CҡU1��Qu��U�ECCU��VEM��]EDb�GVIRC��Q�U�S�B�Q�LA|��p�NFOUN_�DIAG�YRE�X#YZ�cE�WѴh�8�dpqa`T��2�I�M�a�V|be��EGR�ABB��Y�a�LKERj�C4���FC-A�6504x��7u��S BE��h'�`�CKLAS_@l�BA���N@i  G��T$��� @ݲմ$BAƠwj �!q�eb��uTYSp�H����2�šI�t:b�f��B)�E3VE����PK���flx��GI�pNO���2���#�HO����k � ���
8��Pi�S�0ޗ��RO>�ACCEL?0=�-��VR_�U7@�`���2�p��AR��P�A��̎K�D��REwM_But 
�r�JMX �l�t��$SSC�U ����r��QN@m $� �S�P�NS��wLEX�vn T�ENAB 2�W@��oFLDRߨFI�P��t�ߨ(Ğ�?BP}2HFo� ���V
Q MV_PI��8T@󐉰�F@�Z�+�#���8�8#��GA�B���LOO��J�CBx��w"SCON<(P�PLANۀ�Dp�3F�d�v�9PէAM��Q ;����SM0 E�ɥ�8ɥWb72�$`<�8T��,`RK<h"ǁVANC�����R_Ou N@p (��-#<#c��c2_�ACw�A/�N@q 4������`	�^�o�r hn���1^�N&OFF`|�p�`X��`�DEA�
�P�,`SK�DMP6VI=E��2q w��@|���rs < {����4���r{7��D����6�CUSTz�U��t $G��TIT1$P9R\��OPTap �O�VSF�йsu�p��0`r&�@AS�MOwvI�|�ĄJ,�����eQ_WB��	wI���� @O3�@o�XVRxxmr���T���ZA{BC��y op����)�
� �ZD�$�CSCH��z Lu����`�2�%PC ��7PGN ��<�<�A��_FUNH��@	 �ZIPw�{I��LV,SL���~� 
�Z/MPCF��|��E�����X�DMY_L�NH�=�C�� ��}� $�A� ]�CWMCM� C,SC&!���P�� $J���DQ���� ���������_�Q,2�����UX�a\�UXEUL��a�������(�:�(�J���FT�FL��w�C�Z��~Zp+�6�mp��Y@Dp � 8 $R�PU<��> EIGH����#?(�iֱ�b���et� �a����У$B�0�0@�	�_�SHIFD3-�RV2V`Fcв�	$5��C�0��&!�������b
�sx�uD�T�R��V̲��SP9H���!� ,���������4A�RY�P��%������%���"�%!  *�H�(UN0�� �"�2�����K��q0GSPDak����P� �O����0�ĳ���"!NGV�ER`q i�w+I_AIR�PURGE  i  i/�F`�E�Tb�4��)  �� h2ISOLC  �,�"�!�Л!��%��P+�_/*O�B��Dm�?@��!H771  34n?�?�9� �`�E/#�)x� S2;32�� 1i� LTEk@? PENDA�34�1 1D3<�*? Main�tenance /Cons B�? F�"O,DNo UseMJOOnO�O�Op�O�O2�2NPO;�/" 19%�1CH�=� �-Q		�9Q_!UD1�:___RSMAVgAILn�/%�>A!SR  �+���H�_�P1�TVAL�.&���P(.�YV�L�}� 2i��� D?�P 	 �/_oUQNo�orci�o �g�o�o�o�o�o *,>tb��� ������:�(� ^�L���p�������܏ ʏ ��$��H�6�X� ~�l�����Ɵ���؟ �����D�2�h�V��� z��������ԯ
��� .��R�@�b�d�v��� ��п�������(��N�<�r�i�$SA�F_DO_PUL�S. jQp����C�A� �/%�&0S�CR ��`X�����е��4�1IAIE���b  vo$�6�H�Z�l�~�߀�ߴ����������HS��2%��0�d%�@�rb��� @�"k�}���T��h� J`���_ @��T7 ������#�0�T D��0�Y�k�}������� ��������1C�Ugy�O�Ef������  =�5;�o��� 1p�U�
�t��Di�������
?  � ��*�� ����gy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?OO%O7O<A���`OrO �O�O�O�O�O�O�O?O �_._@_R_d_v_�_@�_�_�_�Q _�R0M JTo!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏJO��'� 9�K�]�o�������_ ɟ۟����#�5�G� Y��_�U�_�ҙ����� ϯ����)�;�M� _�m���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������π��0�B�T�f�;� �?�q߮��������� ��,�>�P�b�t�� ������������\����Y���	12345�6781h!B�!����F������������� ���� ��;M _q������ �%7I[l *������� //1/C/U/g/y/�/ �/�/n��/�/	?? -???Q?c?u?�?�?�? �?�?�?�?O�/)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ O_�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�op_�o�o�o /ASew�� �������o+� =�O�a�s��������� ͏ߏ���'�9�K� ]����������ɟ۟ ����#�5�G�Y�k� }���������s�կ��w���0�L��CH  Bpw� �  �=�2��� } �=�
���  	�o�ί��ǿٿ���	r������@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� ��%Ϻ��������� &�8�J�\�n���� �����������"�Q��*�����;�<M����D���  ��]�w�*�Z򛱛�t  d�����*��`*��$SCR_�GRP 1�*P3� �� �*� �6�	 �
�� <�+*�'UC|@�g�y�yD� �W�!�y�	�M-10iA/7�L 123456�7890��� 8��MT� � �#
�	L��	Č� N
���Y���y�
M_	P����� ,?��H�
 ���1/@A/g/y/H�ߙ!T/�/P/�/p3��+���/B�S�!�,?*2C4&Ad�R?�  @s�j5N?�7?���7&2R��?}:&F?@ F�`�2�? �/�?�?OO-OSO>O wObO�O=j1�2�O�O�O�O�DB��O�O;_ &___J_�_n_�_�_�_ �_�_o�_%o�5j�eSgxo6���uo�ox�b�1j16�&J�o�h0�4j9j9B� w��$Y̯@HtA!�Nhcu�/�%pp�	drsq ����zq�x� �� (&�*�2�D�V�o�z�e�������ECL�VL  �����iqpQ@��L_DEFAULT~ ��s��փHOTSTR��qq��MIPOW�ERF��H����WFDO� ��RVENT �1ɁɁ� L�!DUM_EI�P�����j!AF_INE‧���O!FT}�֞��r��!-/� ���F�!RPC_M'AING�)��5���NY�VISb�t�����ޯ!TPѠPU�կ��dͯ*�!
P�MON_PROX	Y+���e�v��D��fe�¿!RD�M_SRVÿ��g���!R,*ϑ�Yh��Z�!
[�M���iIϦ�!RL�SYNC����8|����!ROS|����4��>�!
C}E�MTCOM?߲��k-ߊ�!	S�C'ONS�ߒ�ly����!S�WASRCdݿ��m��"�!S�'USB#n�n�!STMC��o]�����ѳ�����,���P�V�ICE�_KL ?%d�� (%SVCPGRG1S�����2��D����3������4��D����5��6;@��7ch�����9����%�� ������0���� X�����-��� U���}��� / ���H/���p/�� �/��F�/��n�/�� �?��8?���`? ��/�?��6/�?��^/ �?��/X�j��q��� #OhO��lO�O{O�O�O �O�O�O�O _2__V_ A_z_e_�_�_�_�_�_ �_�_oo@o+odoOo �o�o�o�o�o�o�o �o*<`K�o �������&� �J�5�n�Y���}����ȏ���^�_DEV� d��M{C:�4���?GRP 2d�
@��bx 	�/ 
 ,V��o� u�[����������� ٟ���:�L�3�p�W� ������ʯ��� �W� $�ۯH�Z�A�~�e��� ����ؿ�������2� �V�=�zό�sϰ�� ���ϝ�
���.�@�'� d�K߈ߚ߁߾ߥ��� �������<�#�5�r� �ϖ���������� ��&��J�1�n���g� ��������������" 4��X|�u� �����0 )fM�q��� �;�/�>/%/b/ t/[/�//�/�/�/�/ �/?(??L?3?p?W? i?�?��?�?�? O�? $OOOZOAO~OeO�O �O�O�O�O�O_�O2_ _V_h_�?�_C_�_�_ �_�_�_
ooo@o'o doKo]o�o�o�o�o�o �o�oo_Nr Y������� �&��J�\�C���g�ए����ڏ�d ��	ȏ���5� �Y�D�}���%����������ʑv�ʕڟ �ҟ���,��P�^� ����ƙF�����ԯ¯ ����.�p�U���� ��v�����п���6� \�-�l��`�Nτ�r� �ϖ������2ϼ�&� ��6�\�J߀�nߤ��� ��
ߔ�����"��2� X�F�|�ߣ���l��� ��������.�T��� {���D����������� ��\�AS
, t�����4 X�L:\^p� ���0�$// H/6/X/Z/l/�/��/ /�/�/�/ ??D?2? T?�/�/�?�/z?�?�? �?�?O
O@O�?gO�? 0O�O,O�O�O�O�O�O _ZO?_~O_r_`_�_ �_�_�_�_�_2_oV_ �_Jo8ono\o�o�o�o �o
o�o.o�o"F 4jX��o��~ �z���B�0�f� ����V�����Џҏ ���>���e���.� ��������̟Ο��� X�=�|��p�^����� ����ȯ�D��T�� H�6�l�Z���~����� ۿ���Ϡ��D�2� h�Vό�ο���|��� ��
����@�.�dߦ� ����T߾߬������ ���<�~�c��,�� ���������D�)� ;������\������� �����@���4" DFX�|���� ��0@B T����z�� /�,//</���/ �b/�/�/�/�/?�/ (?j/O?�/?�??�? �?�?�?�? OB?'Of? �?ZOHO~OlO�O�O�O �OO�O>O�O2_ _V_ D_z_h_�_�_�O�__ �_
o�_.ooRo@ovo �_�o�ofo�obo�o �o*N�ou�o> �������&� hM�����n����� ����ȏ��@�%�d�� X�F�|�j�������� ,���<�֟0��T�B� x�f���ޟï����� ���,��P�>�t��� ��گd�ο����� (��Lώ�sϲ�<Ϧ� ���ϸ�������$�f� Kߊ��~�lߢߐ��� ����,��#������� D�z�h�������� (���
�,�.�@�v� d������� ������� (*<r��� ��b���� $z�q�J�� ����/R7/v  /j/�z/�/�/�/�/ �/*/?N/�/B?0?f? T?v?�?�?�??�?&? �?OO>O,ObOPOrO �O�?�O�?�O�O�O_ _:_(_^_�O�_�_N_ p_J_�_�_�_o o6o x_]o�_&o�o~o�o�o �o�o�oPo5to�o hV�z���� (�L�@�.�d�R� ��v������$��� ��<�*�`�N���Ə ���t�ޟp���� 8�&�\�����L��� ��گȯ����4�v� [���$���|�����ֿ Ŀ��N�3�r���f� Tϊ�xϮϜ������ ����Ͼ�,�b�P߆� tߪ�����ߚ���� ��(�^�L���ߩ� ��r����� ����� $�Z������J����� ��������b���Y ��2�z���� �:^�R�b �v����6 �*//N/</^/�/r/ �/��//�/?�/&? ?J?8?Z?�?�/�?�/ p?�?�?�?�?"OOFO �?mOO6OXO2O�O�O �O�O�O_`OE_�O_ x_f_�_�_�_�_�_�_ 8_o\_�_Po>otobo �o�o�o�oo�o4o�o (L:p^��o �o�� ��$�� H�6�l�����\�Ə X�֏��� ��D��� k���4�������ҟ ����^�C����v� d���������ί��6� �Z��N�<�r�`��� �������󿪿̿�� �J�8�n�\ϒ�Կ�� �������������F� 4�j߬ϑ���Z��߲� ���������B��i� ��2���������� ��J�p�A����t�b� ����������"�F� ��:��Jp^�� ����� 6 $FlZ���� ���/�2/ /B/ h/��/�X/�/�/�/ �/
?�/.?p/U?g?? @??�?�?�?�?�?O H?-Ol?�?`ONOpOrO �O�O�O�O O_DO�O 8_&_\_J_l_n_�_�_ �O�__�_o�_4o"o XoFoho�_�_�o�_�o �o�o�o0T�o {�oD�@��� ��,�nS����� t���������Ώ�F� +�j��^�L���p��� ����ܟ��B�̟6� $�Z�H�~�l����ɯ ۯ��������2� �V��D�z��������$�SERV_MAI�L  ���~ƸOUTPUTո_�@ʴ�RV 2j�  � (r���<�ʴ�SAVE���TO�P10 2� d 毜Ϯ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~����j�n�YPY�ǳFZ�N_CFG j��=��J�~��GRP 2���g� ,B   �A �D;� B} �  B4=ÿRB21I�H7ELL��j�e��)�*�����%RSR����� �&J5G� k������.?�  ��/�>/P/"\/ ��X/z"{ �U'&"2��dh,g-�"EHKw 1S �/ �/�/�/#?L?G?Y?k? �?�?�?�?�?�?�?�?�$OO1OCO?OMM� S�ODFT?OV_ENBմ��e��"OW_REG�_UI�OȲIMI_OFWDL~@�N��BWAIT�B �)��V��F�YwTIM�E��G_�VA԰_�A_UNcIT�C~Ve�LC�@WTRY�Ge�ʰ�MON_ALIA�S ?e�I%�he��oo&o8oFj�_ io{o�o�oJo�o�o�o �o�o/ASew "������� �+�=��N�s����� ��T�͏ߏ����� 9�K�]�o���,����� ɟ۟ퟘ��#�5�G� �k�}�������^�ׯ �����ʯC�U�g� y���6�����ӿ忐� ���-�?�Q���uχ� �ϫϽ�h������� )���M�_�q߃ߕ�@� �������ߚ��%�7� I�[�������� r������!�3���W� i�{���8��������� ����/ASe �����|� +=�as�� B����/�'/ 9/K/]/o//�/�/�/ �/�/�/�/?#?5?�/ F?k?}?�?�?L?�?�? �?�?O�?1OCOUOgO yO$O�O�O�O�O�O�O 	__-_?_�Oc_u_�_ �_�_V_�_�_�_oo�c�$SMON_�DEFPROG �&���Aa� &*S?YSTEM*obg� $JO0dR�ECALL ?}~Ai ( �}bo@�o�o�o�o�o �o ,>Pbt�� ������(�:� L�^�p��������ʏ ܏� ���$�6�H�Z� l�~������Ɵ؟� ���� �2�D�V�h�z� �����¯ԯ����� �.�@�R�d�v���� ����п���ϙ�*� <�N�`�rτ�ϨϺ� ������ߕ�&�8�J� \�n߀�ߤ߶����� ���ߑ�"�4�F�X�j� |������������ ���0�B�T�f�x�� �������������� ,>Pbt�� �����(: L^p���� �� /�$/6/H/Z/ l/~//�/�/�/�/�/ �/�/ ?2?D?V?h?z? ?�?�?�?�?�?�?�? O.O@OROdOvO�OO��O�O�O�O�O_�@)�copy mc:�diocfgsv�.io md:=�>10.109.�3.62:200A8	_W_i_{_�K3R�frs:orde�rfil.dat� virt:\t/emp\4[6BP�_��_�_o�A+�V*.d�_�[�_Zolo~o�X�
xyzrate 61 (o:oLo�oH�o�U�g�o �o �o]o��U6�_�X?mpback�oO���� }-Sdb%`*�*~�]�o�l���U1x�t:\&� ��8�HpQ�����P2��a����N�Џa� s�����3�N�ߟ� ��(�:�̟]�o�������$SNPX_�ASG 2�������7  R�%���Я�  ?���PAR�AM ��^�� �	��PӤ��PӨ$�������OFT_KB_CFG  ӣ�����OPIN_S_IM  ����}���������RV�NORDY_DO�  )�U���QSTP_DSBi���ϐ�SR }�� � &#��D�O�O�:�TOP_ON_ERRʿ���o�PTN z�����A���RING_PRM�y�ܲVCNT_GOP 2��!���x 	���ϗP��#���Gߔ�VD��RP' 1��"�8Ѩ� *߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�}�z����� ����������
C @Rdv���� ��	*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?[?X?j?|?�? �?�?�?�?�?�?!OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLoso po�o�o�o�o�o�o�o  96HZl~ ��������� �2�D�V�`�PRG�_COUNTJ�9��{�ENB��}��M��L���_UPD� 1'�T  
k�����"�K�F� X�j���������۟֟ ���#��0�B�k�f� x���������ү���� ��C�>�P�b����� ����ӿο���� (�:�c�^�pςϫϦ� �������� ��;�6� H�Z߃�~ߐߢ����� ������ �2�[�V� h�z���������� ��
�3�.�@�R�{�v� ������������ *SN`r����t�_INFO {1�Ҁ� 	 ��3��,B�@-���?!��c΁8:$�p��� D���DH�  C4  ´����YSDEBSUG����� dՉ��SP_PASSB?+LOG� ���  �� ��  ��с�UD1:�\;$�<"_MPC A-셽/�/�x!�/� 쁝&SAV �D)���d!|"�%��(SV�+TEM�_TIME 1:D'�� 0�/�?��.TMEMBK  �сd d/�?��?�<X|Ҁ�3 @�?C�O:O�JLOmOzI�J
! �@p?�O�O�O�C �_ _2_D_V_h_��n_�_�_�_�_�_�_�_o"o\�e1oVoho zo�o�o�o�o�o�o�o 
.@Rdv���O5SK�0�8��`�?���F=� Q4�O%O΄AJ�0[Da YO��}O�M!��O�я�����O!�� �!�t�9�p9�g�y���_L����ӟ���	��� $�C�7og� y���������ӯ��� 	��-�?�Q�c�u���𙿫����T1SV�GUNSPD%% �'%��2MO�DE_LIM �a9"ܴ2�	�� D-۵ASK_OPTION �9!�F�_DI EN�B  U�%f�B�C2_GRP 2A!�u#o?SG��C�����ԼBCCFG 3#��*< ��`ߐI�4�Y� �jߣߎ��߲����� ����E�0�i�T�� x������������/��S�>�w����� t���u�����c��� 	B-f�.��4[  �������  02Dzh�� �����/
/@/ ./d/R/�/v/�/�/�/ �/�(���/?&?8?J? �/n?\?~?�?�?�?�? �?�?O�?4O"OXOFO hOjO|O�O�O�O�O�O �O__._T_B_x_f_ �_�_�_�_�_�_�_o o>o�/Voho�o�o�o (o�o�o�o�o(: Lp^���� ���� �6�$�Z� H�~�l�������؏Ə ��� ��0�2�D�z� h���To��ȟ���
� ��.��>�d�R����� ��z�Я������� (�*�<�r�`������� ��޿̿���8�&� \�Jπ�nϐϒϤ��� ���ϴ��(�F�X�j� �ώ�|ߞ��߲����� ���0��T�B�x�f� ������������� �>�,�N�t�b����� ������������: (^�v���� H���$HZ l:�~���� ���2/ /V/D/z/ h/�/�/�/�/�/�/�/ ?
?@?.?P?R?d?�? �?�?t�?�?OO*O �?NO<O^O�OrO�O�O �O�O�O�O__8_&_ H_J_\_�_�_�_�_�_ �_�_�_o4o"oXoFo |ojo�o�o�o�o�o�o �o�?6Hfx� �������v�&��$TBCSG_GRP 2$�u��  ��&� 
 ?�  Q�c�M���q��� �����ˏ��*�1��&8�d, ��F�?&�	 HCA{��>�ffb��N��CS�B�pI�����V��33��fn�C
��ԝB������&h��Belt�\ԟ�A��!L��;���.�C{��9��������G�w�CHd��k�Ư��C�����@��I�� -���
�X�u�@�R����̻�����	V�3.00I�	mt7���*� �%���ֶ:�H?j� &�H�� N�� �O�  ����a� ϏϘ�*�J21��'8��Ϥ�CFG� )�uB� ,E������d�#��#�I�W��pW� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ��������I�cp "4��gRw�� ����	-? �cN�r��&� �����/</*/ `/N/�/r/�/�/�/�/ �/?�/&??J?8?Z? \?n?�?�?�?�?�?�? O�? OFO4OjOXO�O �O`�O�OtO�O_�O 0__T_B_x_f_�_�_ �_�_�_�_�_�_,oo Poboto�o@o�o�o�o �o�o�o�o(L: p^������ �� �6�$�F�H�Z� ��~�����؏Ə��� �2��OJ�\�n���� ����������
� @�R�d�v�4������� ��ί����ү(�N� <�r�`���������ʿ ̿޿��8�&�\�J� ��nϐ϶Ϥ������� ��"��2�4�F�|�j� �ߎ����߀��� �� ��B�0�f�T��x�� �����������>� ,�b�P���������v� ������:(^ L�p�����  �$H6lZ |������/ �/ /2/h/�߀/�/ �/N/�/�/�/
?�/.? ?R?@?v?�?�?�?j? �?�?�?�?O*O<ONO OO�OrO�O�O�O�O �O�O _&__J_8_n_ \_�_�_�_�_�_�_�_ o�_4o"oXoFoho�o |o�o�o�o�o�o�/ $6�/�oxf�� ������,�>� ��t�b�������Ώ ��򏬏��&�(�:� p�^���������ܟʟ �� �6�$�Z�H�~� l�������دƯ���  ��D�2�T�z�h��� Jȿڿ������
� @�.�d�Rψ�vϬϾ� ���Ϡ������*� `�r߄ߖ�Pߺߨ��� �������&�\�J� ��n���������� ��"��F�4�j�X�z� |������������� 0B�Zl~(� ������, Pbt�D���8���   #� &0/"�$�TBJOP_GR�P 2*���  ?��&	H"O#,V,����x�� =k%  �< �� =�$ @ g"	 �CA��&��SC��_%�g!�"!G��"Q빅�/� .{2^��R=�C�S�?��?��&0L��B�  �B<�'??J7�/�/?�(��6}? ?({�à5;��v 6��*?<?�;B��7C��  D�!�,0ã�B�0OK:��Z�Bl  @p�B@�ff?��
�CH�0��?gO  A�zG�2jG�&�5�333�O�K;�ي|A�!@J@�ffC�Z0zjO�Oz@ǰ��U�O�$#��
0R�E1_CV;xC�sQ@��@&?ff@��O�_ptF�X_�$:�H�R�J=q�_�8AP:��t-�Q?�33@�@@�Oo�_,i$o ZGLo6oDoro�o~o8o �o�o�o�o3�o�RlVd��V4��&b x�%	V�3.00m#mt	7A@�s*�l$!��'� E��q�E���E�]\�E�HFP=�F�{F*Hf�F@D�FW�3�Fp?F�M�F���F�M�F��F�ş�F��F�=�F���G��G.8�CW��RD3l)D���E"��Ex��
E��E�,�)FdRFBF�HFn� F����F��MF����F�,
Gl�Gg!G)��G=��GS5��GiĈ;M@;W�o�|# 2 EdXz&/��&"�?��PYOWOE#�ESTPARS c (a E#HRw�ABLE 1-V)' @�#R�7�Q � �R�R�R��'#!R�	R�
R��R���!R�R�:R���RDI��`!��ԟ���
�r�Oz���������̯ޮ��Sx�^# <����� ÿտ�����/�A� S�e�wωϛϭϿ��� ����;-w�{�_"��6� �1�C�U���%�7��I�[����NUM [ �`!� �$  ��m���_CFG .���B�H IMEBF_T�T}���^#��G�VE�Rk�H�]�G�R {1/�� 8��" �� �A�  ������������  �2�D�V�h�z����� ��������/
e @Rhv���� ���*<N `r������ '///]/8/J/`/n/@�/�/�/�/r���_���t�@~�t�MI_�CHANS� ~� ~!3DBGLVLS��~�s�$0ETHE�RAD ?��
w0�"��/�/�?�?�l�$0ROUTq��!�!�4�?�<SNMASKl8~�}1255.2E�s0O�BOTO�st�OOLO_FS_DI}��%�V9ORQCTRL� 0���#��MT �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo&l�OIo8omoq��PE_DETAI�J8�JPGL_CONFIG 6��ᄀ/cel�l/$CID$/grp1qo�o�o/壀�?Zl~ ���C����  �2��V�h�z����� ��?�Q����
��.� @�Ϗd�v��������� M������*�<�˟ ݟr���������̯@�}a���&�8�J�\���^o��c��`���˿ ݿ���Z�7�I�[� m�ϑ� ϵ������� ���!߰�E�W�i�{� �ߟ�.���������� ��A�S�e�w��� ��<���������+� ��O�a�s�������8� ������'9�� ]o����F� ��#5�Yk�}�����`��User Vi�ew �i}}12�34567890 �//,/>/P/X$� ,�cx/���2�U �/�/�/�/??s/�/�3�/b?t?�?�?�?�??�?�.4Q?O(O�:OLO^OpO�?�O�.5 O�O�O�O __$_�OE_�.6�O~_�_�_�_ �_�_7_�_�.7m_2o DoVohozo�o�_�o�.8!o�o�o
.@��oagr lCamera� �o����� �ޢE�*�<�N��h�z�`�������I  �v �)��$�6�H�Z�l� ���������؟���� �2�Y��vP9ɟ ~�������Ưد��� � �k�D�V�h�z��� ��E�W�I5�����  �2�D��h�zό�׿ ����������
߱�W� ދ��X�j�|ߎߠ߲� Y�������E��0�B� T�f�x�߁ulY��� ������
����@�R� d�������������� ��W� iy�.@Rd v�/����� *<N��W��i �������� /*/</�`/r/�/�/�/�/as9F/�/? ?1?C?U?�f?�?�? D/�?�?�?�?	OO-O
�j	�u0�?hOzO�O �O�O�Oi?�O�O
_�? ._@_R_d_v_�_/OAO �p�{,_�_�_oo)o ;o�O_oqo�o�_�o�o �o�o�o�_�u���o M_q���No� ��:�%�7�I�[� m�NEa����ˏݏ ����7�I�[��� �������ǟٟ���� ͻp�%�7�I�[�m�� &�����ǯ����� !�3�E�쟒�9�ܯ�� ����ǿٿ뿒��!� 3�~�W�i�{ύϟϱ� X�����H����!�3� E�W���{ߍߟ����������������  ��L�^�p���������� ��   "�*�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</�N/`/r/�/�  
���(  �@�( 	 �/�/�/�/ �/? ?6?$?F?H?Z?@�?~?�?�?�?�*2� �l�O/OAO�� eOwO�O�O�O�O��O �O�O_TO1_C_U_g_ y_�_�O�_�_�__�_ 	oo-o?oQo�_uo�o �o�_�o�o�o�o ^opoM_q�o�� ����6�%�7� ~[�m��������� ُ���D�!�3�E�W� i�{�ԏ��ß՟� ����/�A�S���w� ����⟿�ѯ���� �`�=�O�a������� ����Ϳ߿&�8��'� 9π�]�oρϓϥϷ� ��������F�#�5�G� Y�k�}��ϡ߳���� ������1�C�ߜ� y������������� 	��b�?�Q�c���� ����������(� )p�M_q������0@ �������� ��#�frh:\tpg�l\robots�\m10ia4_?7l.xml�X j|�������.��/1/C/U/ g/y/�/�/�/�/�/�/ �//?-???Q?c?u? �?�?�?�?�?�?�?
? O)O;OMO_OqO�O�O �O�O�O�O�OO _%_ 7_I_[_m__�_�_�_ �_�_�__�_!o3oEo Woio{o�o�o�o�o�o �o�_�o/ASe w�������o ��+�=�O�a�s����������͏ߏ��I �<<w  ?�� 4��,�N�|�b����� ��ʟ�Ο���0�� 8�f�L�~���������������(�$T�PGL_OUTP�UT 9����;� $�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ�����$�����2345678901��� � 2�D�V�^����υߗ� �߻�����w����'�9�K�]���}g��� ������o����1� C�U�g���u������� ����}���-?Q c������� ��);M_q 	������ �%/7/I/[/m/// �/�/�/�/�/�/�/? 3?E?W?i?{??%?�? �?�?�?�?O�?OAO SOeOwO�O!O�O�O�O��O�O_�O� $$Ӣ��OW=_o_ a_�_�_�_�_�_�_�_ �_#ooGo9oko]o�o �o�o�o�o�o�o�oC5g}��� �����}@���"�� ( 	 iW�E�{�i����� Ï��ӏՏ���A� /�e�S���w������� �џ���+��;�=��O���s����Ƹ  <<\ޯ� )�ͯ�)��M�_��� ʯ����<���ؿ��Ŀ � �~�$�V��Bό� ��x�����2ϼ�
ߤ� ��@�R�,�v߈���p� ����j�������<� �߬�r������ �����`�&�8���$� n�H�Z���������� ����"4Xj�� R��L���� |Tf �� v��0B//� &/P/*/</�/�/��/ �/h/�/??�/:?L? �/4?�??n?�?�?�? �? O^?�?6OHO�?lO ~OXO�O�OO$O�O�O �O_2___h_z_�O �_�_J_�_�_�_�_o�.o��)WGL1�.XML�cm�$�TPOFF_LI�M Š�p��{�qfN_SVy`�  �t�jP_�MON :����d�p�p2miS�TRTCHK �;���f~tbVT?COMPAT�h*q��fVWVAR �<�mMx�d R e�p�bua�_DEFPROG7 %�i%|��rd_DISPLA�Y�`�n�rINST�_MSK  �|� �zINUSE9R �tLCK)��{�QUICKMEN�M��tSCREl����+rtps�c�t)������b��_桉STz�iRAC�E_CFG =��iMt�`	nt
�?��HNL 2!>�z���T{ zr@� R�d�v���������К��ITEM 2?�,� �%$12�34567890<�%�  =<�C�<U�]�  !c�k�wp'���ns�ѯ5� ���k������j�ů ��鯕���A�1�C�U� o�y�󿝿I�oρ�� ��	��-ϧ�Q���#� 5ߙ�A߽�����e߳� �����M���q߃�L� ��g��ߋ����%� w� �[���+�Q�c� ��o��������3��� {�;������G _����/�Se .�I�m�� �=�a/3/ ������k// �/�/�/]/?�/�/�/ ?�/u?�?�??�?5? G?Y?�?+O�?OOaO�? mO�?�?�OO�OCO_ _yO+_�O�Ox_�O�_ �O�_�_�_?_�_c_u_ �_o�_Wo}o�o�_�o o)o;o�o�oqo1C �oO�o�o��% ��[��Z���S�@��_�� 3 ے_� ����y
 Ï�Џ�~��UD1:\����q�R_GRP� 1A �� 	 @�pe�w�a�@��������ߟ͞�� ��ّ�>�)�b�M�?�  }���y��� ��ӯ������	�� Q�?�u�c���������Ϳ�	-���o��SCB 2B{� h�e�wωϛϭ���������e�UTORIAL C{���@�j�V_CON?FIG D{��������O�OUTP�UT E{�����������%� 7�I�[�m����� ���������%�7� I�[�m���������� ������!3EW i{������� �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/��/??'? 9?K?]?o?�?�?�?�? �?�/�?�?O#O5OGO YOkO}O�O�O�O�O�O �?�O__1_C_U_g_ y_�_�_�_�_�_�O�_ 	oo-o?oQocouo�o �o�o�o�o�_�o );M_q��� ���yߋ����-� ?�Q�c�u��������� Ϗ���o�)�;�M� _�q���������˟ݟ � ��%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ���
�� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� ��������������� 1CUgy�� �����	- ?Qcu��������/�x���$/6/ !/a/� �/�/�/�/�/�/�/? ?'?9?K?]?�?�? �?�?�?�?�?�?O#O 5OGOYOkO|?�O�O�O �O�O�O�O__1_C_ U_g_xO�_�_�_�_�_ �_�_	oo-o?oQoco t_�o�o�o�o�o�o�o );M_q�o �������� %�7�I�[�m�~���� ��Ǐُ����!�3� E�W�i�z�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�π�'�9�K�]�o�~���$TX_SCRE�EN 1F8%w  �}�~�@��������
���� m&��\�n߀ߒߤ߶� -�?������"�4�F� ��j��ߎ������� ��_����0�B�T�f� x������������� ��>��bt� ���3�W (:L^���� ����e/�6/�H/Z/l/~/�//�/��$UALRM_M_SG ?����� �/���/�/)?? M?@?q?d?v?�?�?�?�?�?�?O�%SEV7  �-EF�"ECFG H�Ż��  ��@�  AuA   ;Bȁ�
 O�� �ŨO�O�O�O�O__�&_8_J_\_jWQAGR�P 2I[K 0���	 �O�_� I�_BBL_NOT�E J[JT��l�������g@�RDEFPR�O� %�+ (% O.o��oUo@oyodo �o�o�o�o�o�o�o�?�\FKEYD?ATA 1K�ɞP�p jG�� h_���P����u,(J����J� 1�n�U�������ȏ�� ����"�	�F�X�?� |�c�������֟�������0��T��~�� d���������ӯ寈� y�� �2�D�V�h��� ������¿Կ�u�
� �.�@�R�d�v�Ϛ� �Ͼ������σ��*� <�N�`�r�ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |�������������� ��0BTfx� ����� �>Pbt��o� ����//:/ L/^/p/�/�/�/5/�/ �/�/ ??$?�/H?Z? l?~?�?�?1?�?�?�? �?O O2O�?VOhOzO �O�O�O?O�O�O�O
_ _._�OR_d_v_�_�_ �_�_M_�_�_oo*o <o�_`oro�o�o�o�o Io�o�o&8J �on�����W ���"�4�F��j��|�������ď֏��܋�������)��K�]�7�,I���A�����֟� ϟ��0�B�)�f�M� �������������ݯ ��>�%�b�t�[��� ���ο����(� :�L�[�pςϔϦϸ� ����k� ��$�6�H� Z���~ߐߢߴ����� g���� �2�D�V�h� �ߌ���������u� 
��.�@�R�d���� �������������� *<N`r�� ����&8 J\n���� ����"/4/F/X/ j/|//�/�/�/�/�/ �/?�0?B?T?f?x? �?�/�?�?�?�?�?O O�?>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_�_5_ �_�_�_ oo$o�_Ho Zolo~o�o�o1o�o�o �o�o 2�oVh z���?��� 
��.��R�d�v��� ������M����� *�<�ˏ`�r������� ��I�ޟ���&�8��J�!0L��!0���u�����q���ͯ��,������"� 	�F�X�?�|�c����� ��ֿ������0�� T�f�Mϊ�qϮϕ��� �������,�>�?b� t߆ߘߪ߼�˟���� ��(�:�L���p�� ������Y��� �� $�6�H���l�~����� ������g��� 2 DV��z���� �c�
.@R d������� q//*/</N/`/� �/�/�/�/�/�/�// ?&?8?J?\?n?�/�? �?�?�?�?�?{?O"O 4OFOXOjO|OSߠO�O �O�O�O�OO_0_B_ T_f_x_�__�_�_�_ �_�_o�_,o>oPobo to�oo�o�o�o�o�o �o:L^p� �#���� �� �6�H�Z�l�~����� 1�Ə؏���� ��� D�V�h�z�����-� ԟ���
��.���R� d�v�������;�Я� ����*���N�`�r�����������@��}��@����@��	��+�=��,)� n�!ߒ�y϶��ϯ��� ���"�	�F�-�j�|� cߠ߇����߽����� ��B�T�;�x�_�� ��O��������,� ;�P�b�t��������� K�����(:�� ^p����G� � $6H�l ~����U�� / /2/D/�h/z/�/ �/�/�/�/c/�/
?? .?@?R?�/v?�?�?�? �?�?_?�?OO*O<O NO`O�?�O�O�O�O�O �OmO__&_8_J_\_ �O�_�_�_�_�_�_�_ ��o"o4oFoXojoq_ �o�o�o�o�o�o�o�o 0BTfx� �������,� >�P�b�t�������� Ώ������(�:�L� ^�p��������ʟܟ � ����6�H�Z�l� ~������Ưد��� ���2�D�V�h�z��� ��-�¿Կ���
�� ��@�R�d�vψϚ�)� ����������*�`�,��`���U�g�y�Qߛ߭���,���ߑ����&� 8��\�C���y�� �����������4�F� -�j�Q���u������� �����_BTf x�������� ,�Pbt� ��9���// (/�L/^/p/�/�/�/ �/G/�/�/ ??$?6? �/Z?l?~?�?�?�?C? �?�?�?O O2ODO�? hOzO�O�O�O�OQO�O �O
__._@_�Od_v_ �_�_�_�_�___�_o o*o<oNo�_ro�o�o �o�o�o[o�o& 8J\3���� ���o��"�4�F� X�j��������ď֏ �w���0�B�T�f� ����������ҟ��� ���,�>�P�b�t�� ������ί�򯁯� (�:�L�^�p������ ��ʿܿ� Ϗ�$�6� H�Z�l�~�Ϣϴ��� ������ߝ�2�D�V� h�zߌ�߰������� ��
��.�@�R�d�v�h���qp���qp���������������,	N� r�Y������������� ��&J\C� g������� "4X?|�m �����/�0/ B/T/f/x/�/�/+/�/ �/�/�/??�/>?P? b?t?�?�?'?�?�?�? �?OO(O�?LO^OpO �O�O�O5O�O�O�O _ _$_�OH_Z_l_~_�_ �_�_C_�_�_�_o o 2o�_Vohozo�o�o�o ?o�o�o�o
.@ �odv����M ����*�<��`� r���������̏��� ��&�8�J�Q�n��� ������ȟڟi���� "�4�F�X��|����� ��į֯e�����0� B�T�f����������� ҿ�s���,�>�P� b��ϘϪϼ����� �ρ��(�:�L�^�p� �ϔߦ߸�������}� �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z�	�����@��������
��������5GY1{�g, y�q��� <#`rY�}� ����/&//J/ 1/n/U/�/�/�/�/�/ �/�/ݏ"?4?F?X?j? |?���?�?�?�?�?�? O�?0OBOTOfOxO�O O�O�O�O�O�O_�O ,_>_P_b_t_�_�_'_ �_�_�_�_oo�_:o Lo^opo�o�o#o�o�o �o�o $�oHZ l~��1��� �� ��D�V�h�z� ������?�ԏ���
� �.���R�d�v����� ��;�П�����*� <�?`�r��������� ��ޯ���&�8�J� ٯn���������ȿW� ����"�4�F�տj� |ώϠϲ�����e��� ��0�B�T���xߊ� �߮�����a����� ,�>�P�b��߆��� ������o���(�:� L�^������������ ����}�$6HZ l�������� y 2DVhz�Q�|�Q�����������,�/./�/R/9/ v/�/o/�/�/�/�/�/ ?�/*?<?#?`?G?�? �?}?�?�?�?�?OO �?8OO\OnOM��O�O �O�O�O�O�_"_4_ F_X_j_|__�_�_�_ �_�_�_�_o0oBoTo foxoo�o�o�o�o�o �o�o,>Pbt ������� �(�:�L�^�p����� #���ʏ܏� ���� 6�H�Z�l�~������ Ɵ؟���� ���D� V�h�z�����-�¯ԯ ���
����@�R�d� v��������Oп��� ��*�1�N�`�rτ� �ϨϺ�I������� &�8���\�n߀ߒߤ� ��E��������"�4� F���j�|������ S�������0�B��� f�x�����������a� ��,>P��t �����]� (:L^��� ����k //$/ 6/H/Z/�~/�/�/�/��/�/�/���+�>�����?'? 9=?[?m?G6,YO�? QO�?�?�?�?�?OO @ORO9OvO]O�O�O�O �O�O�O_�O*__N_ 5_r_�_k_�_�_�_�_ ��oo&o8oJo\ok/ �o�o�o�o�o�o�o{o "4FXj�o� �����w�� 0�B�T�f�x������ ��ҏ������,�>� P�b�t��������Ο ������(�:�L�^� p��������ʯܯ�  ���$�6�H�Z�l�~� �����ƿؿ���� ��2�D�V�h�zό�� ����������
���_ @�R�d�v߈ߚߡϾ� ��������*��N� `�r����7����� ����&���J�\�n� ��������E������� "4��Xj|� ��A��� 0B�fx��� �O��//,/>/ �b/t/�/�/�/�/�/ ]/�/??(?:?L?�/ p?�?�?�?�?�?Y?�?� OO$O6OHOZO�$�UI_INUSE�R  ����{A� � [O_O_MENHIST 1L{E�  �( �@��)/�SOFTPART�/GENLINK�?current�=menupag�e,1133,1`�O_ _2_�?� �O�M936�O�_�_�_ �_TR�_�_ oo$o6o Ho�_lo~o�o�o�o�o Uo�o�o 2D�o hz�����c �
��.�@�R��v�@��������Џ���o� �Ao���0�B�T�f� i���������ҟ�s� ��,�>�P�b��� ������ί�򯁯� (�:�L�^�p������� ��ʿܿ�}���$�6� H�Z�l�~�Ϣϴ��� ���������2�D�V� h�zߌߏϰ������� ��
��.�@�R�d�v� ���)��������� ���<�N�`�r����� %���������& ��J\n���3 ����"�� Xj|����� ��//0/�T/f/ x/�/�/�/�/O/�/�/ ??,?>?�/b?t?�? �?�?�?K?�?�?OO (O:OLO�?pO�O�O�O �O�OYO�O __$_6_ H_3E~_�_�_�_�_ �_�O�_o o2oDoVo �_�_�o�o�o�o�o�o uo
.@Rd�o ������q� �*�<�N�`�r���� ����̏ޏ����&��8�J�\�n�Y_��$�UI_PANED�ATA 1N������  	�}��ǟٟ0����!� )#�G� cT��r���������̯ 3��ׯ�&��J�1� n�U�������ȿ���p���"�\Y� kQG�Z�_�qσϕϧ� �����P����%�7� I�[�m��ϑ�xߵߜ� ���������3�E�,�i�P������6� �榓���*�<�N� `�����Ϩ������� ��i�&8\C ��y����� �4Xj���� ������M/ ��B/T/f/x/�/�/�/ /�/�/�/�/?,?? P?7?t?�?m?�?�?�? �?�?Ow�:OLO^O pO�O�O�?�O�O=/�O  __$_6_H_�Ol_S_ �_�_�_�_�_�_�_�_  ooDoVo=ozoao�o O#O�O�o�o
. @�od�O���� ��I���<�#� `�r�Y���}�����ޏ ��׏���8�J��o�o ��������ȟڟ-��� q"�4�F�X�j�|��� ������֯������ 0��T�f�M���q��� �����W�i��,�>� P�b�t�ǿ�Ϫ���� ������(ߏ�L�3� p߂�iߦߍ�������  ���$�6��Z�A�~���}������������"�)��G���6� s�����������4��� ����K2oV ���������#�����$UI�_POSTYPE�  �� 	 /�U�QUICKMEN  ds�W�RESTORE �1O� � ��� /#���m+/T/f/ x/�/�/?/�/�/�/�/ ?�/,?>?P?b?t?/ �?�?�??�?�?OO (O�?LO^OpO�O�O�O IO�O�O�O __�?_ 1_C_�O~_�_�_�_�_ i_�_�_o o2o�_Vo hozo�o�oI_So�o�o Ao�o.@Rd �����s�� �*�<��oI�[�m�� ����̏ޏ�����&� 8�J�\�n��������xȟڟ�SCRE��?�u1�sc�u2�3��4�5�6�7r�8��TAT`�� ��MUS#ER�����T���Sks���4��5���6��7��8��UN�DO_CFG aPd����UPDX�����No�ne���_INF�O 1Q�<��0%��W���E��� i���������տ� ��:�L�/�pς�eϦ���)�OFFSET' Td@���{� �����	��-�Z�Q� cߐ߇ߙ��ϝ����� �� ��)�V�M�_�q� �۹�����
����t��)�WORK U4�����A�S���ψ�UFRAME�  ���&�RTOL_ABRT���$���ENB����G�RP 1V��?Cz  A� ��+=Oas������U������MSK  �<���mN��%4��%��<)��_EVN������>�2W��
� h��UEV���!td:\e�vent_use3r\-�C7���}�F��SP���spotwel=d�!C6����!�Z/�/ :'�H/~/l/�/�/�/ �/-?�/Q?�/? ?�? D?�?h?z?�?O�?)O �?�?OqO`O�O@ORO �OvO�O_�O�O7_�O�[__Z]W+�2X�����8V_�_�_  �_�_o�_,o>oobo toOo�o�o�o�o�o�o �o:L'p��]����$VA�RS_CONFI��Y�� FP{����|CCRG��\��>�{�t�D.� BH� pk�a��C�� ��}�?�x��C,&Q=��ͩ��A �MR2bN���	}�	���@�%1: SC�130EF2 *(����{�����X� ˂5}�����A@vk�C�F� w�Q�[���|�����������T����\��ϟ �\� B���;�e�@�ǟ`��� ��S�����̯���ۯ �&�}��\�G�Y���pE���ȿ�TCC�Ac
��������p�GF�pgd���-�23456789017�?��ׁ$���4�v�Nm�� ��϶�BW�����i�~}�:�o=LA� څ�6�@�6�ͿZ���$i�7����(��W��� -�]�X�jĈߚߕϳ� ����������%�7� I�r�m�ߨ�ߵ��� �������8�3�E�W� ������}��������� ����/�A�S�e�w��MODE��t ��RSLT e�|k�%"zς�� ;�1��d��`�>�SELEC���c��	IA_WO֗Pf �� }W,		���|���G�P ������RTSYNC�SE� ��$�	#W�INURL ?*ـ�;\/n/�/�/�/�/�uISIONTMOU���A#� ��%�gSۿ��SۥP��� FR:\�#\�DATA\�/ ��� MC6L�OG?   U�D16EX@?\�'� B@ ���2T1���?�?�?\������� n6  ���GV�2\�� -��5�� �  ��Z�@U0>58TRAINj?��4*B{Rd_Cp��F'#`{2�'$�":��h#� (�kI �Mw��O�O�O�O�O1_ _U_C_]_g_y_�_�_\�_�(STA� i�B�@�?o0o�:$o\bo�%_GE�j#�;�~@ �
�\�|�btgHOMIN�_kSۮ��`�2(,,��CWǖBve�JMPERR 2=l#�
  Qo�: ��"�4Fwj| ��������l�&%S_g0RE鰹m�^۴LEXdn��1-ehoVM�PHASE  �e׃BޱOFF� _ENB  ޢ$VP2�$oS�ۯ��x�c C�;�@ �@�;���?Gs33'D*AA���]� ��0ޱ�`r}�XC��܅���\A8-۟E ���� ��#�5��������� ����}��������� �c�X���A�����ϯ �+��߿��M�B� q���xϊϹ���Ϸ� ������7�I�;�m�b� )ߣ�Eߓߡ߳���� �3���W�L�{ߍ��� �����������/� $�6�e�W���c�y��� �����������O� ��?M_q����� ��'9�=7 Is������ /m/%/3/E/s��TD_FILTE:�`s�k �x2�`����/�/�/�/�/ 	??-???Q?�6�/~? �?�?�?�?�?�?�?O� OoiSHIFTM�ENU 1t}<5�%5�~O)�\O�O �O�O�O�O�O�O'_�O _6_o_F_X_�_|_�_��_�_	LIVE�/SNAP�Sv�sfliv���_�{z`ION ҀyU
`bmenu&o�+o�_�o�oV"<E�uZz��4IMO�v����zq�WAITD�INEND  0�ec��b�fOKو'OUT�hSDywTIMdu��o|G�}#�{C�zbx�z�xRELE���ڋxTM�{�d��c_ACT`و���x_DATA 	wz���%�oď5Fx��RDIS
`E��o$XVR�ax�n��$ZABC_G�RP 1yz�.�� ,�2̏.M{ZD��CSCH�`�z���aP@�h@6�IP�b{'����şן�[�MPC�F_G 1|'����0�r�8��� �}�'��p�s� �	(���  <�l0  ��?���������D��ƣH�1w�쯛�����ѯ F���m!#��{��@�ܵ�� /�C4  ´ſ׾ĸ� �	��1�?�i���'��0�����	��`�~����_CYLI�ND~!� ��� ,(  * .�?ݧ+�h�Oߌ�s� ��������(�	� x�-��&�c�߇�� ������j�P����)���~�_�q��� �2�'��� �&���� ������&��I��cA���SPH�ERE 2��� �������A� T/A��e�� ����/N` =/�a/H/Z/�/��/��/�/�ZZ� � �f