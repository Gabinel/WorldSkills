��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� � P�COUPLE,  o $�!PPV1GCES C G1�!��PR0�2	 � $SOFT��T_IDBTOT_AL_EQ� Q1�]@NO`BU SPI�_INDE]uEX�BSCREEN_��4BSIG�0�O%KW@PK_F�I0	$TH{KY�GPANEhD� � DUMMYE1d�D�!U4 Q�!RG1R�
 � $TIT1 d ��� 7Td7T� 7TTP7T55V65V75V85V95W05W>W�A�7URWQ7UfW1pW1
zW1�W1�W 6P!�SBN_CF�!-�0$!J� ; |
2�1_CMNT�$FLAGS]n�CHE"$Nb�_OPT�3�(C�ELLSETUP�  `�0HO��0 PRZ1%{cM�ACRO�bREP	R�hD0D+t@��bl{�eHM MN�yB
1�UTOB �U�0 �9DEVIC4ST	I�0�� P@13�r�`BQdf"VAL�#ISP_UNI��#p_DOv7IyFR_F�@K%D13�x;A�c�C_WA?t��a�zOFF_@N.�DEL�xLF0q8�A�qr?q�pF�C?�`�A�E�C#��s�ATB�t�d��MO� �sE �� [M�s��2�R;EV�BILF��1�XI� %�R � � OD}`j�_$NO`M� +��b�x�/�"u��� ����!X�@D�d p E R�D_Eb��$F�SSB�&W`KBD�_SE2uAG� G
�2 "_��B�� V�t:5`ׁQC �a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR�B�IGALLOW�� (KD2�2�@VAR5�d!�AB �e`BL[@S � !,KJqM�H`S�pZ@�M_O]z����CFd X�0G�R@��M�NF�LI���;@UIR�E�84�"� SWIYT=$/0_No`S�"�CFd0M� =�#PEED��!��%`���p3`J3tV�&$E�..p`L�>�ELBOF� ��m��m�p/0��CP�� F�B����1���r@1J1E_y_T>!Բ�`��g����G� �0WARNMxp�d�%`��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqM��� R�r$ORIأ.&ӧRT�SF\g CHGV0I�Ep�T��PA�I{��T�!��� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5��6�7�8�9��4��x@�2 @.� TRQ��$%f��4ր����_U����z��Oc <� �����Ȩ3�2��LL�ECM�-�MULTIV4�"$��A
2q�CHILD>�
1���z@T_1b  4� STY2�b4�=@�)24����@��� |9$��T��A�I`�E��eTOt���E��EXT����ᗑ�B��22(�0>��@��1b�.'��}!�A�K�  �"K�/%�a��R���N?s  =�O�!M���;A�֗�M�� 	��  =�I�" �L�0[�� R�pA��$JOBB�����ނ�TRIGI�# dӀ����R�-'r0��A�ҧ��_M��b7$ tӀFL6�BsNG�A��TBA�  ϑ�!��
/1�À�0���R0�P/p ����%�|��Bqh@W�
2JW�_RH��CZJZ�_zJ
?�D/5C�	�ӧ�t�@��Rd&�������ȯ�qGӨg@N�HANC��$LG /��a2qӐ� ـ@��!A�p� ���aR��0>$x��?#DB�?#3RA�c?#AZt@�(p.�����`FCT��ƕ�_F࠳`�SM��!I�+lA�%` � ` ���$/�/����[�a��M�0\��`l��أHK��AEs@�͐�!�"W��N� SbXYZW�`�"�����6	��I���'  . I�I��2�(p�STD�_C�t�1Q��US�TڒU�)#�0U�[�%?IO1��� _Up�q�* \��=�#AORzs8Bp�;�]��`O6  RSY�G�0�q^EUp��H`�G�� ��]�DBPX�WORK�+* $SKP_�p��A��TR�p , �=�`����Z m�O1D3��a _C"�;b�C� �GPL:c�a�tDőS�D�W�3B�b����P�.� &)DB�!�-�B APR��
I�Ja3��. /�u������K�LuY/�_�����0�_���PC��1�_���~�EG�]� 2�_�SVP�RE.��R3H �$C��.$L�8c/$uSނz IkI3NE�WA_D1%�ROyp�������q0�c7 t@�fPA���?RETURN�b��MMR"U��I�C�Rg`EWM@�SIGNZ�A ��|�e� 0$P'��1$P� m�2�p�p'tm�+pD��@ �'�bdNa)r�GO_AW ��@4ؑB1I�CSd�(�KCYI�4���`1w��qu��t2�z2�vN��}��E}sDEV�Is` 5 P �$��RB��I�wPk��I_BYȧ��"�T7Q�tHN{DG�Q6 H4���1�w��$DSBLC��o��vg@��|tL��7O�f@]���3FB���FEra8��ׂ�t}s���8> pi�T1?���MCS����fD �ւ[2H� W ��EE���%F����t����9 T�p��x�NK_N:�����UZ��L�wHA�vZ' ~�2���P~r�q7w: �=MDLn��9�ጂٱh����! e����J��~� +����,�N�D����3���ՒG!aqSL�Ad�7;  ��INP��"�����}q_ V�4<�06`C� �NU��  D�L�ק��SH!�7=BM��q���ܢӢ����g���>P +$ٰ�٢��^��^�Y�FI B�\��Ă��'A	'AW�l�NTV��]�V\~�X�SKI�#T� ��a�ۺ�T1J�3:39_�P�SAFN����_SV�EXCSLU��N@�DV@�Ll @�Y����S�H�I_V
0\2PPL5YPRo�HIM�T��n�_MLX��pVORFY_�Cl�M��gIOC�UC_� �����O�q�LS(�0v�FT4Q���)��@P�E$�t��A��CNFt�6եup��pm�4ACHD��o������AFC C	PlV�TQTP?�� ί� ?`�@TA��@�0L@ ��N���]� @����T��T! S����te@{R�A DO�� w23���!n��	_1�#�H!�̔�΀�K��B�2��MAR�GI�$���A ���_SGNE�C;
$�`�a^aR0 ��3��@ B��B��ANNUN�P?����uCN@�`%0��`��� ���BEFc@]I�RD @Q�F���4OT�`�sFTӠHR,Q��CQ0�M��N�I|RE�����A�W���DAY=CLOCAD�t;T|�<S5}�EFF_AXI��%F`1QO3O��Eq���@_RTRQ�E�G����0RQ
�2Evp ��|��F�0f�R0 �tM��AMP�E<� H 0�`œ^��`Ds�DU�`��v�BCAr� I?��`N ErIDLE_PWRI\V!n0�V�wV_[ |�� ��DIAG�5J�o 1$V�`SE�3TQl�e��P�l�^E_��Y�VE6� �0SWH�q (� �b|�Gn�3OHxPPHZ�IRAl�B�@�[� �a�b�1�w3�O  � ��v�|�I�0 ��pRQDW�MS-�%AX{6Y�LIFE�@�&�MQy�NH!Q%��F#�C����CB0�mpNr$�Y @�aFLAl�f��OV0]&HE��>l�SUPPO�@u��y��@_�$��!_�X83�$gq�'Z�*W��*B1�'T�#`�k2XYZáY�Y2D8CY`T@�`N�����f� �C�I2��IC�TA�K `�pCACH�ӫ�3�����I��bNӰUFFI� \��@��;T��r<S6CQ.�MSW�5�L 8	�KEYI7MAG�cTMLa���*Ax�&E���B��OC�VIER-aM ���BGL����y�?G� 	��П4N�m:�ST�!�B P�D,P�D��D��@�EMAI䐔a��M��r�FAUL|RO bB�c�� spUʰMA�"`T'`E�P< �$S�S[ � ITw�BUF�7y��7r�tN[�LSUB1T��Cx�o�R�tRSAV|U>R'c2�\�WT���P�T�*`S�n�_1PbU���YOT(�bK��P��M��d����WAX��2��XX1P��S_GH#
���YN_���Q <�Q�D��0���M��� T�F�`�|�\�DI��EDT�_Pɰ:�R��b�G�RQM�&��Jq�a����׀��Fs� S (�SVqpB��4��_�.��a��T�� �@���B�SC_R]1IK>B'r��$t�R"A#u�H�aDS�P:FrP�lyIM@|Sas�qz��a� U>wh� <1%sM�@IP��0s��0`tTHb0ЃdTr��T`asHS�c�CsBSCʴq0� V`�����S�_D��/CONVE�G���Hb0^v1PFHy�dCs�`&a?ASC���s�MERg��aFBC�MPg��`ET[� �UBFU� DU�%P�D�:12�CD�Wy�p�P�CG�[@N	O6�:�V� ��� �R��P���C������w��A��`��W/H *�LƠ�C c�W����Y�賂��� ��q�|���A*��7}�8}�9}�H T���1��1��1��U1��1ʚ1ך1䚕1�2��2����2���2��2��2ʚ2�ך2�2�3��3R��3����3��3��U3ʚ3ך3�3�94��QEXT[�X[b�H``t&``z�k`t˷$���FDR�/YTPV��RpK"	��K"REM*9F��]"OVM:s/ŽA8�TROV8�D�T�PX�MXg�INp8ɉ W��INDv�BH2
�ȕ`K ^`G1a �a��@Q%7Da��RIV��u"]"GE[AR:qIO.K(�H4N�`���,(�F@|� I3Z_MCM<0.K! �F� UT����Z ,�TQ?� b�y@t�G?t�E |�.�>Q�����[ �Pa�� RI�E��UP?2_ \ �@=S#TD	p<TT����p�����a>RBACUbG] T��>R�d)�j�%C�E��0��IFI���0��i�{�4�PT�T��FLUI�D�^ �?0gHPUR �gQ�"�r�a�4P�+ I�$��Sd�k?x��J�`CO�P��SVRT��N�x$�SHO* ��CAS�S��Qw%�pٴBG_%��3���<�FORC�B��^o�DATA��_�BKFU_�1�bb�2�a�m=mm�b0��` �|��NAV	`)������$�S�Bu#?$VISI���2SC	dSE������V��O�$&�B�K�� ��$PO���I��FM�R2��a  ��	��`#��@&�8�O� (�_��9��+IT_^�ۄ�)M�����DGC{LF�DGDY�LD����5Y&��Q$RY�M됇CbN@{	? T�FS�P�D�c P��W�cK �$EX_WnW1P%`]��"X3�5�s�G+�d ���ָ�SWeUO�DE�BUG��-�GRt��;@U�BKU���O1R� _ P�O_ )�����M���LOOc>!SM E�R�a��u _E� e >@�G_�TERM`%fi'��ORI�ae gi%y�SM_�`>Re !hi%V�(ii%3�UP\Bj� -����e��w#� f���G�*ELTOr�A�bF�FIG�2��a_���@�$�$g$wUFR�b$�01R0օ� OT_7F��TA�p q3NST��`PAT�q�0�2P'THJ�ԀE�@�c3ART�P'58�Q�B�aREL�:�aSHFT�r�a�1�8E_��R��у�& � 	$�'@i�
����sN@bSHI�0�Uy�= �QAYLO�p� Oaq�����1����pERV��XA��H�� m7�`�2%�P�E3�P��RC���ASYM�a��aWJ07����AE�ӷ1�I��ׁUT@�`Oa�5�F�5P�sXu@J�7FOR�`M # �O!k]��`5&�0L0��`HOL ;l �s2T�����OC1!E��$OP��qn����$�����$��PR�^��aOU��3e���R�5e�X�1 �eo$PWR��IMe�BR_�S�4�� �3��aUD��k�Q�dm���$H�e!�`AWDDR˶HR!G�20�a�a�apRR��[�n H��S����%���e3��e���e��SE���z�HS�MNu�o���Pªq��0OL�s߰`ڵ<�I ACRO��&1��ND_C�s��A<fdK�ROUP��R!_�В� �Q1|�= �s���y%��y-��x�� �y���y>�=A�����AVED�w-��uy&sp $�І�P_D�� ��'rP�RM_���!HT�TP_�H[�q (ÀOBJ��b �[$˶LE~3��>\�r � ����J��_��TE#ԂS�P�IC��KRLPiHI�TCOU�!��L ���PԂ������PR���PSSB�{�JQUERY_FLAvs��@_WEBSOC����HW�#1��s��`<PINCPU(���O���g������d��t��O� �IwOLN�t 8��yR��$SL!�$INPUT_�U!$`��P �G֐SL.���u���2�.��C��B��IOa�F_AS:=v�$L+ਇ+�A��bb41�����Z@HYʷ�����#qe�UOP:w `v�ϡ˶�¡�������"`PIC`����� �	�H�IP_ME���v�x Xv�IP�`(�R�_N�p�d����Rʳp�ױQrSaP �z�C��BG(��� ��M�Av�y lLv@CTApB��AL TI�3UfP_ ۵�0�PSڶBU_ ID � 
�L � `�Q0��L��0z)�����ϴ�NN�_ O��I�RCA_CNf� �{ �Ɖ-�CYpEA������� �IC�ǫ�tpR�=Q�DAY_
��NTVA�����!��5�����SCAj@��CL��
����
���v�|`5�VĬ2b�l�N_�PACV�n�
���w�})� T��S�����
��e����T� 2| Ր�� �v�~��֣�ذLAB1��_ �חUNIX��ӑ ITY裪��e~�p�� ���<)���R_U�RL���$A;qEAN ���s`vsTeqwT_U��m�J��X�M�$���E��"��R祪�� A�,�2��JH���FLy���= 
���
�UJ]R|U� ���F��6G��K7��D>�$�J7�s��J8*�7����3�E�7��&�8�\�)�APHI�Q4�y�DkJ7Jy8R��L_KE'�  �K͐L}MX� � <U��XRi�����WATCH_VAZqu@Aស�FIEL`��cy�n���:� � u1VbwPCTX�j��Y �LGE���� !��LG_SIZ΄�[8Zm�ZFDeIYp1! gXb ZW �S`� 8�m��� �b ���A�0_i0_CM c3#�*'FQ1�KW d(V(Bbpo pm�p� |Io�1 pb p�W RS��0  M(C�LN�R�۠-�DE6E3��� �c�i���PL#�7DAU"%EAq�͐�T8". GH�R��y��BOO�a��3 C��F�ITV�l$�A0��RE���(SCRX����D&�ǒ�qMARGI�Sp�,@����T�"�y�S���x�W�$y�$��JG=M7MNCHt�y�FN��6K@7r�>9�UFL87@L8FWDvL8HL�9STPL:�VL8"�L8s L8RS"�9HOPh;��C9D�3 R��}P�'IUh�`4@�'�5$ ��S2G09�pPOWG�:�%�3,�64��N9EX��TUI>5I� �ӌ���� �C3�C<0'�,�o�:��&�@�!NaqvcAcNAy��Q�AI]�8gt7Ӝ�DCS���c�RS�cRROXXOdWS��ÂRoXS{X�(IGNp 
Ђ=10 ��[T�DEV�7LL���CZ!*�C �	 8�Tr$f/蛒����Z�3A�a�	 W�h萦�Oqs�S1Je2Je3Ja��BSPC G� �ƋG`-T� �%��Q�T�r@�&E�V�fST�R9 YBr~�a �$E�fC�k�g��f	v��CB� L����� �� u�xs뀔�g�q�jt:��!�#_ ����ʐv�#Ӡ �s �M�C�� ���C�LDP᠜�TRQ�LI ���y�tFL ���rQ��s5�D���w�~�LD�u�t�uOR�G���1�RESERV��M���M�Œ�C�s��� � a	�u�5�t�uSV���p��	1�����RCLMC��M�_�ωxА��: MDBGh��I����$DEBUGMAS������JU�$T8P��EF��d�
�MFRQ~Ҥ� � K	�HRS_RU��bq��A��$EFRE�QUu!$0YOVER�k��f��PU1EFI�%�Gq�� �6�Y�z��� \����E�$U��`��?��
�P)SI`��	��CA ���ʲ�σUY�%�?�( 	��MISC��� d��aRQ���	��TB� � 1���A��AX���|����EXCESg��d�M�H�9��u���9d�SC�` O� H�х�_��@���������pKE�a��+�� &�B_, �FLICBtB� QoUIRE CMOt�QO���r�LdpMD�� �p{!��5b����ND!��I�!���L �D;
$�INAUT�!
$R#SM�ȧPN����C�PSTLHᗻ 4U�LOC�fR�I"��eEX��ANqG.R.���ODA]���q��� �RMF0����icr�@mu8���$�SUPiu��FX��IGG! � ���cs�F� cs
Fct��ޒ�b5��` E��`T�5�tC��g�#TI��7�M���7� t��MD���A)��XP��ԁ��H��.���DIAa��Ӻ�AW�!��0af���D@#�)֡O�㥀��� -�CUp V	����.����!_��� ��{`�c������� |�P|��0� ��P�{�KEB��e-$qB��o�=pND2ւ�����2_TXltXGTRAXS������LO: ����}� ���C�.�&���RR2h���� -�!A�� ?d$CALI����GFQj�2F`RIN�bn�<$Rx�SWq0ۄ���ABC�ȇD_J��{�q��_�J3��
��1SPH, �q�P����3��(H�9pq�#J�34n���O�QIM�M�CSKP�zb7?SbJ+�M�Qb�y8����_AZ��/��EL�Q.ցOC�MP��N�� RTE�� �1�0 ����1��@ ZScMG�0����JG�p�SCLʠ��SPH�_�PM��f��q��u�RTER��n��Pk�_EP�q�`A0� �cM��DI�Q�23UdDF  쀐�LW�VEL��qINxr�@�_BALXP.��Y/�J�0�'$Q�IN���B]�C�9%�".�8!:6p_T� �F%a"�6#a!��k)�Q�DHʠ��\�9`�$Vw��_�A$�=����&A$���S�h��H ��$BEL� m��_oACCE� 	8<�0IRC_�q��@�NT��c$SPSʠ�rL��� M4�s9 .7��GP/6��9�7$3�73S2T�͡_Ga�"�0�1��8�17_MG}�DD�1���FW�p��3�5$3�2�8DEKPPA�BN[7ROgEE �2KaBO�p�Ka���1�$USE_tv�SP��CTRT�Y4@� �� <qYN�g�A�@�FR �ѢAM:�N�=R�0O�v1�DINC(��B�4����GY��ENC�L���.�K12��H0IN¿bIS28U��ONT|�%NT23_���fSLO���|P��Iذ~��V�~�$���hpU#�CQ MVMOSI�1<�[�1��M�PERCH  �S��� �W���SlщR ��l����E�0�0P	AS2EeL�DP7�O�NUЉZ�f�VTRK�RqAY"�?c��a S2�e�c�����BP�MOM�B���C�H�}�Cj��c�3gBT��DUX �2S_BC?KLSH_CS2Fu :��V���C-�esRoz|�A�CLALMJTp@��`� �uCHKe |����GLRTYp� ��8T��5���_�ùT'_UM3��vC3��1�Z���LMT��_ALG��%���0�E*� K�=�)�@5F�@8 9��Nb��)hPC�Q)hHpТ��5�uCMC��\�0�7CN_��N��L�;SF�!iV�B���.W���S2/�ĈCAT�~SH�Å��4  V�q/q/V�T1�f�0PA�t�B_P�u�c_f Z�f�Pe�cݔ�uJG���ѓ��OGއ�TORQU~@�S�i @e��R� @B�_Wu�d@�!a��#`��#`�Ih�Iv�I�#F��S�:X��I�0VC00��֢1ܮ�0�⦇JRKܬ!��<�D�BXMt�<�M�_sDL�!_bGRVg�``��#`��#A�H_%�8?��0��COS��� ��LN#���ߥŴ�  ��=������꼰�<�1Z���VA�MYǱ:���᯻[�THET=0�UNK23�#��l�#ȰCB��CB�#Cz�AS�ѯ����#����SB�#��'GTSkZAC�����&���$DU�phg6�j��E�%eQ%a_��x�NEhs1K�t�� y��A}Ŧկ׍�����LCPH����^U��Sߥ ����������!��(Ʀ�V��V�غ ��UV��V��V
�V�UV&�V4�VB�H��@������d�����H
�UH�H&�H4�HB�O��O��Os���O���O��O
�O�O*&�O4�O(�F�Ҫ��	���SPBA?LANCE_J�6�LE��H_}�SP�>!۶^�^��PFULCb�q����K*1�UTO_<�p�uT1T2�	
22N�q2VP�M�a�� i�Z23	qTu`O��1Q�INSEG2�QREV�PGQgDIF�ep)1�U6�1��`OBK�q�j�w2,�VP�qI�L�CHWAR4B�"A�B��u$MEC�H��J��A��vAX��aPo���׫"� �� 
�?�10UROB�PCRS2#%Ղ����C1_ɒT �� x $WEgIGH�@�`$��d\#��I�A�PIFvAN�0LAG�B��S�B�:�BBIL�%OD��`�Ps"ST0s"P�:�pt �!N�C!L ��P 
P2�Aɑ  �2��Tx&DEBU҄#L|0�"5�MMY9C59N��$4�`g$D|1 a$0�ېl� ���DO_:0AK!� �<_ �&� �q�A��B$�"� NJS�8_�P�@���"O�p �� %�T7P?Q��TL4F0TICK,�#�T1N0%�3=pB�0N�P� u3�PR\p��A��5��5U0PR�OMP�CE�� $IR"��A�p8BX`wBMAIF��A�BQE_� OCX�a��@RU�COD�#F9U�@�&ID_�P�E�82B> G_SUFF�� �#�AXA�2DO�7/�5� �6GR�#��DC�D ��E��E-��DU4� u�_ H_FI�!�9GSORD�! R 236s�HR�A>N0$ZDT�E�P|�!X5�4 *WL_NA�1�0�R�5DEF_I�X�RF �T�5�"�6�$�6�S�5�UFISm�#�m1|Ј�40c�3�T6�44􁆂�"D� ?rfd�#�D�O@ l2LOCKE���C�?OG2a�B�@UM�E�R�D�S �D�U�D>b�B�c�E�S �Dd�B�&2v2a�C� ʑ�E�R�E�S�C9wwu�H�0P} d�0,a�ТF0W�h�u�c� ��TE�qY4� }�!LOMB_�r��w0s"VIS��I�TYs"AۑO�#A�_FRI��~SI,a�n�R�07��0R7�3�#s"W�W��Q��%�_���AEAS{#�B��|�x`WB�8�45�55�6|#ORMULA_I����G�W� h �
>75COEFF_O�1&)��1���Go�{#S� 52CA�� :?L3�!GRm� � � $�`4�v2X�0TM�g��`�e�2�c��3ERIqT�d�TAP�  ��LL�Dp`S��_S�Vkd��$�vAP��.���AP� ��SwETU,cMEAG@��@Πt �!HRL � g� (�  0���l��l��aw��RH�0�a�a}d]�d��B��Ay`Gax`��t[Ѐk@REC[Q:q��1SK_A y��� P_!1_USER����*���VEL�����-�!��IzP� �M�T�1CFG��� � �0]O�NGOREJ �0l���~[�� 4 e�8��"�XYZ<S��� 3� ��_ERRK!� U ѐ�1�@Ac�Ȱ�!�>�B0BUFINDX����p� MORy�� H_ CUȱ�1���dAyQ?�I>Q	$ +�a����� �\�G{�� � $SI�h��@2	��VOv�q�- OBJyE| w�ADJUF2�yĈ�AY�����D��OUKP����AMR=�T��-���X2DIR����X8f�1  DYNt�0�-�T� ��R��0� ~���OPWOR��� �,B0SY�SBU����SOP�o���z�Uy�XP�`K���PA�q��Ӭ���OP�@U����}�"1��IMA�G۱_ �п"IM�.���IN������RGOVRD"ё�	���P����  >gplcC��L�`BŰ?l�PMC_E�P�1EN��Mr�1212�R�"�SL| ��� ��R OVSL=S��rDEX\a`��2�:�_"���P#����P������2�C� �P>���#�_Z�ERl���:����� @��:��O�@R	Iy��
[�g@e����s�P�PL���  $FREEY�EEU�~�Z��L����T�� ATU9Sk�,1C_T�����B������p�Vc18��P��� Dc1������LQ����MQ��ۡL�XE��x�5I�P�W�` ��UP��H`&aPX;@���43�� �PG�Y��g�$SUB����q���JMP�WAIT~ ���L�OW���1wē CV!F_A�0��R�Z��CC �R$��28IGNR_PL��/DBTB� P*a�#BW@.t�U�0-�IG��!@I�TNLN,�RBѡb�yN!@��PEED~ >��HADOW� ��t���E������PwSPD��� L_ �A�нP���	#UN�q � �RP (�L�YwPa����PH�_PK���b�RETRIE��x������� H�0NFI���� ���V �$ 2}�d�DBGLV<?LOGSIZz�baKKTU���$D�n�_TXV�EM�!Cڡ��� �-R�#�r>��CHECKz��(��L���ϰq)ҹL��NPA�`T�J"����)1P����
�AR�"�BC =Sa��O�@����ATT S�u䡳&� w�^a�3�-#UX^�4�PL��@Z�� $d��qS�WITCH�h�W���AS��f�3L�LB��� �$BA�Dvc��BCAMi��6I��(@#J5��N�UB6[F
A_KNOWK3qB"ЍU��AD+Hc� D���IPAYLOAq�9p�C_���GrѼG�Z�CLqAj��PL�CL_6� !@4��BOA?�T7�VFYCӐ�Jp��D��I�HRՐ�G�TBd��6�J��zQ_J�A: �B�AND���`�T�BQ�q��PL@?AL_ ��0 P=�TAe��pC��D�C�E���J3�P�V�{ T�PDCK^��)b��COM�_AL3PH�ScBE<�߁��_�\�X�x\� �� ���OD_�1�J2�DDM�AR�<�h�e�f�cQ�TI�A4�i5�i6��MOM(��c�c�c�c�cV�B� AD�cv�c\v�cPUBP�R�d�<u�c<u�b}"�1���� L$PI$� �pc��G�y��I�yI�{I�{I�s�`�A ���v��v�J�bp��a��HIG�3 ���0���5Ѐ0�f�?�5N�5�SAMPD Ƣ�0���8�;@�S ��с 6���1���� ���` ���`1�K�P��`腽P2�H��IN1��P ��8�T�/��:�z�Q��z���GAMM&�S|��$GET�d����D^d>�
$�P�IBR��I��$HI��_���1���E=��A�9�*�LW�W�N�9�{�*�Zb����QCdCHKh0�j�ݠnI_�� M�JļRoh�Q ��s�J�-v��S ý$�X 1�N�I��RCH_D�$RN���^�LE@��i�p�Zh8�ţ_MSWFL/M�P7SCR�75�Ҽ ��3�"Ķ�6��`��`ع�紙��0SV���P'������G�RO�g�S_SA�=AH�=ńNO^`C i�_d=��no�O�O �x�ʚ��p�B�u�ȐcDO�A��!�ں �*�t�:�Z1f�;�7լ���C etMmu�o � �YL�snQ ��� ���"��<s�	�����nQ�8��<3M_Wl���A��\p��(�o�MC ��P���Q���ȇ�hpM.�pr� !��!��$�WM��ANGL�!�AM�6d K�=dK�DdK��TT7�ANk@��3�#�PXC 	OEc�QZ��hp	nt�� ���OM� ��ϑϣϵ����`� �c�Z0���hp^a_�2� |a�J��i ���c���cJ��j������jA�{ �{����{ �@{�P�1�P�MON_QU�� �� 860QCO�U��QTHxH�O��B HYS�0ESPBB UE- 3�f0]O�4�  c P��^�RUN_TOʹ�gpO��� �P�@��IND9E�#_PGRA���0���2��NE_NO���ITf��o INFO��a"��ژ��H�OI� =(*�SLEQ!�*0�*�Q OS��l4�� 460ENA�By� PTION��3��r��^GC]F�!� @60J�,�Q���R�d!���u�PEDITN�� �� ��KAQj"� �E(�NU'�(AUTY�%CO�PYAQ�2,�qe�M��N< @+��PRU�Tm� C"N�OU��2$G��$
�R�GADJ��u2X_��IX����&���&W�(P�(~��&9�� z
�N�P_CYCy�{w�RGNSc9�{�s�LGO£��NYQ_FREQ�SrW@��X1�4�L��@�2P0�!�c@�"�CcRE��MàIF�q��NA��%�4_}Gf�STATU~�<f��MAIL��|CyIq�=LAST�1�a*4ELEMg�� ��QrFEASIt;�ւΰ��B"� F�AF����I� ���O2�E u�vBAB$��PE� =�VA�FzQ�I��TqU[��R���S�FRMS_TRpC�Qc��C��Z�
��1�D � ,2ns�؆�	MB 2� `���N�3V�R 2WR*���шR^W�wNj�DOU�^�N��,2PR`�h�1G�RID��BAR�S!�TYuBOT�Op�� |_"�4!� �R�TO��d�� � ����P�OR�c~vbSReV�0)"dfDI[�T�`;aNd�pXg
�XgQ4Vi��Xg6Vi7ViI8:a�Fʒg�z ?$VALU�C0��3D1@(1F05��C !pf���S�1�-ȆAN/��b�1R��]11ATOTALX����=sPWE3I�Q>StREGENQzfr��X�H�]5	v( cTR�CS�Qq_S3��wfp�V�!��r��BE�3�PG0B�( nsV_H�PDA(��p�S_Ya���i6�S��AR(�2� }�"IG_SE�3ȿpb�5_� �tC_��V$CMPl��D�Ep�G���IšZ�~�X�
�% Fm�HA{NC.� p Q�r�2���INT�9`cq�F���MAsSK�3�@OVRMP �PD�1-��W� ��aХT�l�_RF|�{�V�PSLGP�
g�9�j5��,��;pDpS���4��1U���|�TE���`G���`k���J^�<Y�y3IL_Mx4�s��p��TQ( ����@����V.�C<�P�_ �R�F�M]�V1V\�V1j�2y�2j�U3y�3j�4y�4j� ��p۲������ܲ;IN�VIB8�6��#��*�2&�22�3*&�32�4&�42���6�|�J�  �T ?$MC_FK `� �L>�J�х1p�Mj�Iу��zS ���1���KEEP�_HNADD��!H鴓@�C��0	��Q����
�O!�v ঱�p
�և
�REM!�	�Cq�RF�]�b��U�4e	�HPWD�  �SBM����PCOLLAB�*�p��/q�2I�T/0��""NO1�F�CALp⎵��� �, �FLv�A$�SYN���M��C�k��RpUP_DL�Y��zDELAh9�Dq�2Y AD(���(0QSKIPNO�� �`� O��cNT����c�P_�  ��׾ ��cp���q�� ���o`��|`�ډ`��@�`�ڣ`�ڰ`��9�!O�J2R0  �lX�@TR3H��1AH��� �H���$ RD�Cq��� � R"�R, 5��R�1��8E��5TRGE�_C��RFLG"���9W�5TSPC�1�UM_H��2TH�2N}Q�;� o1� y�ED�Q>02 � D� ˈ<��@2_PC3W��S���1Y0L10_�Cw2$C+��� � $\� U@ ��V7�����0� �� c�\����� r@d��C�Q,��7���DZ Gs�RUVL1b[�1h���10]�_DS�������PK ;11�� lڰ�0���q��AT?��$ �Q[7�� ��K 5Tx���HOME�S *�c2h�n������]�`3h���!3EW `4h�h@z�����5h���	//-/?/W6h�b/t/�/�/�/��/ ���!7h��/�/??'?9?�8h�\?n?�?�?�?�?� _S����  �Aa{p��3��+�_�Ed� T0=�nD4vnCIO䑎I�I@`�O��_OP��E�C.rfBXPOW=E	�� X@��f��$$C�d�S����_��5�3�3� �@�sSI��GP�0�QIRTU�AL�O
QAAVM_WRK 2 7U� ?0  �5Qn_rzXk_�] �\A	�P�]�_3�8P��_�_�Ve�\#m/o�Q`5ojo|o�dHPBS��� 1Y� <Xo�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯz�bC$�AXLM�@tiAQ��c  d��IN����PRE�
�E�J�-�_U�P��[�7QHPIO�CNV_�� �	�Pr�US>��g�c{IO)�V 1U[P $E`��Qս9lҿ8P?��i@��� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������ );M_q��� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o��o�m�LARMRECOV a���-���LMDG ���ɰ�LM?_IF ��� ை����zv����%�6�, 
 6�_��r漅�������̍$w���׏���8�J�\�n����NGTOL  a�� 	 A   ���ț�PPINFoO ={ <v�����1��   I�3�a�"rP���t��� �����ί���>�o����j�|������� Ŀֿ�����0�B��PzPPLICAT�ION ?����J��Handling�Tool �� �
V9.30P/�04ǐM�
88g340�å�F0����202�ťʚϬ�7DF3��M̎��NoneM�F{RAM� 6���Z�_ACTIVE��b  sï�  ~p�UTOMODz��A���m�CHGAoPONL�� ���OUPLED 1ey� �������g�CUREQ �1	e{  T�
��	p��w����#r���e�HN���{�HTTHKY��
$r��\[�m���� O�	�'�-�?�Q�c�u� ������������ #);M_q�� ����% 7I[m��� /���/!/3/E/ W/i/{/�/�/�/?�/ �/�/??/?A?S?e? w?�?�?�?O�?�?�? OO+O=OOOaOsO�O �O�O_�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_oo#o5o GoYoko}o�o�o�o�o �o�o1CU gy������ �	��-�?�Q�c���1�TO��|�p�DO_CLEAN��|n��NM  �� �B�T�f�x����%�DSPDRY�R��m�HI���@ /�����,�>�P�b��t���������ίj�MAXa�ۄ��������Xۄ������p�PL�UGG��܇�ӌ�P�RC��B� ���ׯF�OK���ȔSEGF��K������ �.�����,�>�v���LAPӟ澨�� �϶����������"��4�F�X�j߯�TOT�AL�7���USE+NUӰ�� �������1�RGDISPWMMC����C��&��@@Ȓ��Oѐ������_STRI�NG 1
��
��M��Sl��
A�_ITEM1K�  nl�g�y�� �����������	�� -�?�Q�c�u����������I/O S�IGNALE��Tryout M�odeL�Inp���Simulat{edP�OutOVERRА� = 100O�In cycl�P�Prog A�borP���S�tatusN�	H�eartbeat�J�MH Fauyl��Aler�	 ������*8<N` ׃G� ׁY�c����� ////A/S/e/w/�/��/�/�/�/�/�/wWOR��G�-1�?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO8�O�O�NPOE� �@E;�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo�BDEV�Nu`�Obo�o �o�o�o�o�o, >Pbt��������PALT ��E?�A�S�e�w� ��������я���� �+�=�O�a�s����GRI�G뽑1��� ���	��-�?�Q�c� u���������ϯ�� ��)�����R�a� ՟;���������ѿ� ����+�=�O�a�s���ϗϩϻ���O�PREG��y���-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_��q����$ARG_�-0D ?	������� � 	$��	+[��]����������SBN_CONGFIG���� ��CII_S?AVE  ��)����TCELLSETUP ���%  OME_I�O����%MOV�_Hn�����REP�d�����UTOBA�CKY���#��FRA:\�� �����)�'`l ���&� 7"�� 24/0�6{  09:35:24�����͓0������@+=Oas�Ƅ �������/ 1/C/U/g/y/�//�/ �/�/�/�/	?�/-???�Q?c?u?�?�?p�� � _��_\AT�BCKCTL.TM���?�?�?O O��INI�Y�-�~��MESSAG9��GA)��RKODE_QDs�<��zHOw`��O��PAUS�@ �!��� , �	�����O�G,		�O__?_)_ ;_u___�_�_�_�_�_��_�_�_)m�D�@TSK  �M&,O���UPDT�@EGd��`�FXWZD_E�NBED��fSTApDE��e��XIS�?UNT 2��&��(�� 	\`�h�� Q�� �Q�`)�3�������q � Cp�Y,t:p�5�p�JUg~q|�P t����E3�����Dm�w�%�G����aMETrc�2LfE� P q�Bb�B�B��B5RB�G�B���CM\���}?yo�?٥�@?��=@u��?z�R@i����}SCRDCFoG 1��' �A�&�������ԏ�����Q =���H�Z�l�~����� 	�Ɵ-����� �2�`D���域���GR�`��`�O���0NA����	��_ED�C@1n�� 
 ��%-�0EDT�-q����%�p�à�u���������������  ��B��2����*�R�b B���*�q���ϧ���3bϮ�@Ͻϯd?���@��=�O���sϏ�4.� ��{�����W���	����?ߏ�5��j�G�� ��#������}�6��6��Z�����Z� ���I��7��� ��&��λ�&m�������8^ҿ���� 	͇�9K�o��!9*�w��	�S���;��CR ����B/T//�/���w//��РNO_�DEL����GE_�UNUSE���I�GALLOW 1���   (�*SYSTEM�*is	$SER�V_GR�;B0�@REGK5$m3i|B0�NUMp:�3�=P�MU� iuLA�Y�pi|PM�PALD@�5CYC10�.�>�0�>CULSU�?�=�2�A�M3LOWDBOX�ORIt5CUR_�D@�=PMCNV6�6D@10�>�@T4DLI�`=O_9�	*PROGRA�J4PG_MI�>�OPAL�E_U�PB7_B>$F�LUI_RESU`�7p_z?�_�TMRY>h0�,�/�b�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv����������"LAL_OUT 1;�l���WD_ABO�R�0?d�ITR_�RTN  �����g�NONSTO�Ǡ�� 8CE_�RIA_I0���ۀ��ŀFCFG ��۔��o_LIMY22ګ� �  � 	i�J��<e�g��5�� 9���������
���u��P}AQPGP 1�����Q�c�u�b4�CK0����C1���9��@���PC��CUV��]��d��l��as��P���C[٤Um��v�������_�� C����-�m��?�ÂHE� �ONFI�Pq�G�G�_P�@1� �%�������ǿٿ�����G�KPAU�SaA1�ۃ  �2�W��Eσ�iϓ� �ϟ����������#߀I�/�m��eߣ��M~��NFO 1"�;�� �7�������B���ƓA�&����ߌ��I�@��8� A  �%Cj��D����3���7�lB� 3�E�ŀ�O�c�COLLECT_�a"�[�����EN�@p��y���k�NDE���"�3�"1�234567890��\1�� ��֕	H&��)M�r�\,L� ^���]+���������� ��C 2�Vh z������ 
c.@R�v����������� ����IO !���q���u/�/ؙ/�/C'TR�2"'-(׀^)
��.R��#R-�*W� 9_MkOR�$� �;� l5��l9�?r?�?�?�?P�;E2��%S=,W�I?@�@��C׀K)D*ցC�R�&u�XO�WAWBC4  A�jq��׀x׀A"@_Cz  B�@CG��B8��AC  @�yB�׀ց:d��43 <#ׁ
�E���I�O�C=AIJ��'GM?�C�(S=��Qd=AT_DEFPROG �;�%�/m_APINU�SE�V�ۅ�TKEY_TBL  s��ہ���	
��� !"#$%�&'()*+,-�./�:;<=>�?@ABCDPGH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������Ga��͓���������������������������������耇����������������������$��PLCKp�\���P�PSTAn���T_AUTO_D�O��NFsINDx���n��R_T1wT2N����5ŀ�TRLCPLETE����z_SCRE�EN ��kcscÂU��MMENU 1)O� <�[_#�q�� ,�a���>�d���t��� ӏ����	�����Q� (�:���^�p������� ̟�ܟ�;��$�q� H�Z����������Ư د%����4�m�D�V� ��z���ٿ��¿�!� ��
�W�.�@ύ�d�v� ���ϬϾ������A� �*�P߉�`�r߿ߖ� ���������=��&� s�J�\������������'�,�p_MA�NUAL�EqDB�
12�v�iDBG_oERRLIP*�{h! 0��������g�NUMLIM�s:QOE�@DBP�XWORK 1+�{��>Pbt���-DBTB_�q �,��kC3!VD�!DB_AWAYzo�h!GCP OBs=��A�_AL���o�k�Y�p�uO@`�]_�� 1-�+@�
-k-6[��_MM+pIS�`�@"@��ONTIM�wM�OD��&
�U�;MOTNEND��_:RECORDw 13�{ ��[CG�O�f!T/[K ��/�/�/�/_(�/�/ f/?�/??Q?c?�/? �??�?,?�?�?OO �?;O�?_O�?�O�O�O �O(O�OLO_pO%_7_ I_[_�O_�O�__�_ �_�_�_l_!o�_,o�_ io{o�o�oo�o2o�o Vo/A�oeP ^�
���R� ��=��a�s���� ����*�ߏN���'� ��ԏ]�̏�������� ɟ۟v���n�#���G��Y�k�}���TOL�ERENC�B��0� L��g�CS�S_CNSTCYW 24	�t���.������0�>� P�b�x���������ο�����(�:�äD�EVICE 25ӫ ��ϟϱ� ����������/�A���ģHNDGD 36ӫ� CzT�.!�ơLS 27t� S�����������/��U�ŢPARAM 8Gb�A�ՔտRBT 2:�8�<���C�kA� ·���  � A����.SB���A�B��  ���0������.��  X����A�A�C��`��c�u����C�A�CD��k�pz�YA�A��HA�c�� A�	�?(uL^�p���A�Bt/{�D��C��_� 	 A=���ABffA#33�AҊ���A�,A�Cf��a��A��J��7B]���B��Bff�Bᴠ�33C$0.@R� (�� ��A����
/� �//)/;/�/_/q/ �/�/�/�/�/�/�/<? ?%?r?I?[?m??�? �?�?�?�?&O8O�PO bOMO�OqO�O�O�O�O �O_�OOL_#_5_ �_Y_k_�_�_�_�_ o �_�_6oooloCoUo go�o�o�o�o�o�o  �o	h�O�w� ����
��.�	_ _I'�1_�q����� ���ˏݏ���%� r�I�[���������� ǟٟ&����\�3�E� W����ȯ���ׯ� "��F�1�j�E�s��� ��m�������ѿ�0� ��f�=�O�a�sυ� ���ϻ�������� '�9�Kߘ�o߁����� [����(��L�7�p� ��m��������� ��$�����l�C�U� ��y�����������  ��	V-?�cu ����
��@ +dO�s��� �����*///`/ 7/I/[/m//�/�/�/ �/?�/�/?!?3?E? �?i?{?�?�?�?�?�? �?�?FO�jOUOgO�O �O�O�O�O�O__� 'O9OO=_O_�_s_�_ �_�_�_�_�_�_oPo 'o9o�o]ooo�o�o�o �o�o�o:#5 ��O����� ���$��H�Fz�$D�CSS_SLAV�E ;����w��`�_�4D  w���A�R_MENU <w� >�؏���� �2�^rǏ\�n�\����SHOW 2=>w� � fr[q ����Ə�����,� >�D�b�t��� ���� ҟϯ����)�P� M�_�q���������˿ ݿ���:�7�I�[� ��|Ϧ��ϵ������� ��$�!�3�E�l�fߐ� �ߟ߱��������� �/�V�P�z�w��� �����������@� :�d�a�s��������� ��\���*�H�N�K ]o������� �28�GYk }������ "�1/C/U/g/y/�/ ��/�/�/��//? -???Q?c?u?�/�?�? �?�/�??OO)O;O MO_O�?�O�O�O�?�O �?�O__%_7_I_pO m__�_�O�_�O�_�_ �_o!o3oZ_Woio{o �_�o�_�o�o�o�o Do-Se�o��o ������.��=�O���CFG �>�����q��d�MC:\��L�%04d.CSV�\��pc�������A- ՃCH݀z�v�Pw�#��q����:�J�8�7���JPQ�j�)�́�p+��n�RC_OUT [?z������a�_C_FSI �?�� |�����@�;� M�_���������Я˯ ݯ���%�7�`�[� m��������ǿ�� ���8�3�E�Wπ�{� �ϟ����������� �/�X�S�e�wߠߛ� �߿��������0�+� =�O�x�s������ �������'�P�K� ]�o������������� ����(#5Gpk }����� � HCUg�� ������ // -/?/h/c/u/�/�/�/ �/�/�/�/??@?;? M?_?�?�?�?�?�?�? �?�?OO%O7O`O[O mOO�O�O�O�O�O�O �O_8_3_E_W_�_{_ �_�_�_�_�_�_oo o/oXoSoeowo�o�o �o�o�o�o�o0+ =Oxs���� �����'�P�K� ]�o�����������ۏ ���(�#�5�G�p�k� }�������şן ��� ��H�C�U�g����� ����دӯ��� �� -�?�h�c�u������� ��Ͽ�����@�;� M�_ψσϕϧ����� ������%�7�`�[� m�ߨߣߵ������� ���8�3�E�W��{� ������������� �/�X�S�e�w����� ����������0+ =Oxs���� ��'PK ]o������ ��(/#/5/G/p/k/ }/�/�/�/�/�/ ?�/�??H?C?U3�$D�CS_C_FSO ?����1� P [?U?�?�?�?�?�? O
OO.OWOROdOvO �O�O�O�O�O�O�O_ /_*_<_N_w_r_�_�_ �_�_�_�_ooo&o OoJo\ono�o�o�o�o �o�o�o�o'"4F oj|����� ����G�B�T�f� ��������׏ҏ��� ��,�>�g�b�t��� ������Ο����� ?�:�L�^����������ϯʯܯg?C_RPI~>�?�;�d�_� 
�}?.�p����ݿj>SL�@���9�b� ]�oρϪϥϷ����� �����:�5�G�Y߂� }ߏߡ���������� ��1�Z�U�g�y�� �����������	�2� -�?�Q�z�u������� ������
)R M_q����� ��*%7Ir m�����/ �ϛ�,�/W/�/{/ �/�/�/�/�/�/?? ?/?X?S?e?w?�?�? �?�?�?�?�?O0O+O =OOOxOsO�O�O�O�O �O�O___'_P_K_ ]_o_�_�_�_�_�_�_ �_�_(o#o5oGopoko }o�o�o�o�o�o �o HCUg�� ������ �����NOCODE �@������PRE_CHKg B��3�A 3���< ��7��������� 	 <�����?#ۏ%�7� �[�m�G�Y������� ٟ�ş�!����W� i�C�����y�ïկˏ ������A�S�-�_� ��c�u���ѿ����� ��=��)�sυ�_� �ϻϕ��������'� 9���E�o�I�[ߥ߷� ����������#���� Y�k�E���{���� ��������C�U�� =�����w��������� 	����?Q+u� a������ );_qg�Y� �S����%/� /[/m/G/�/�/}/�/ �/�/�/?!?�/E?W? 1?c?�?���?�?o? �?O�?�?AOSO-OwO �OcO�O�O�O�O�O_ �O+_=__I_s_M___ �_�_�_�_�_�?�_'o 9oo]oooIo�o�oo �o�o�o�o#�oG Y3E��{�� ���o�C�U�� y���e����������� 	��-�?��K�u�O� a���������͟�� )��1�_�q��}��� ����ݯ�ɯ�%��� 1�[�5�G�����}�ǿ ٿ�������E�W� 1�{ύ�G�u����ϯ� �����/�A��-�w� ��c߭߿ߙ������� ��+�=��a�s�M�� ��ϑ�������'� �3�]�7�I������ ������������G Y3}�i���� ����C/ y�e����� ��-/?//c/u/O/ �/�/�/�/�/�/�/? )?�?_?q?K?�?�? �?�?�?�?�?O%O�? IO[O5OO�OkO}O�O �O�O�O_�O3_E_;? -_{_�_'_�_�_�_�_ �_�_�_/oAooeowo Qo�o�o�o�o�o�o�o +7aW_i_� �C�����'� �K�]�7�i���m�� ɏۏ�������G� !�3�}���i���ş ������1�C��g� y�S�e���������� ѯ�-���c�u�O� ������Ͽ�ןɿ� )�ÿM�_�9�kϕ�o� �����Ϸ������ I�#�5�ߑ�kߵ��� ��������3�E��� Q�{�U�g������� �����/�	��e�w� Q��������������� +Oa�I� ������ K]7��m� ����/�5/G/ !/k/}/se/�/�/_/ �/�/�/?1???g? y?S?�?�?�?�?�?�? �?O-OOQOcO=OoO �O�/�/�O�O{O�O_ �O_M___9_�_�_o_ �_�_�_�_oo�_7o Io#oUooYoko�o�o �o�o�o�O�o3E i{U����� ���/�	�S�e�?� Q�������я㏽�� ��O�a������� q���͟������� 9�K�%�W���[�m��� ɯ�����ٯ�5�+� =�k�}���������� ���տ�1��=�g� A�Sϝϯω����Ͽ��������Q�c�����$DCS_SG�N CS�����#M�25�-JUL-24 �09:54 E��06��N��39������� X�L��������������ДќM��?Þ�j������{�VERSION� ��V4�.2.10�EF�LOGIC 1D�S��  	D���X�k�X��z�M�PROG_E_NB  ��b���Л�ULSE  ����M�_AC�CLIM��������WRSTgJNT����w�EMO���ѷ�L��INIT EZ��O��OPT_S�L ?	S�1�
 	R575��V��74��6��7��)5A��1��2��l����G�h�TO  �t���.H�V?�DE�X��d����FP�ATH A��A�\4���HC�P_CLNTID� ?+�b� �l�����IAG_�GRP 2JS�� ��a[�D�  D��� D  B߫  B�@ff��/B�@[���W�@�q���B�N�C�-�Bz��Bp@�e`��mp3�m7 7890123456�*�[���  Ao��mAj1Ad�A]�
AW|��AP�AJ-�AC/A;�ǞA4H���@�W  A��A�A3!�_A�@@��B4�� ��t����
�uƨApf�fAj�yAeK��A_�AY���AS� MC�AF��A@ �O��+/=/O$O�c K�w(@�X?8��@��y�/�/�/�/��/8�;d�2�5�?@~ff@x1�'@q��@kC��@d�D@]��@Vv�6?H?Z?�l?~?8s�0l���@e@^���@W\)@O���@H�0?<@7K�@.V�?�?�?�?|
O8S@M00�G<@A��@<�1@5��@/l�@(Ĝ@!�0�\NO`OrO�O�O x'g�L_K�;_�_�__ g_�_�_�_�_o�_�_ �_YokoIo�o�o+o�oX�"� 2�17A�@�J>��R
q?��33?Y��r{��J7'Ŭ2q�63p4�F>r�{�LJ@�p�Zr��
=@�@��Q�jq��@G A�h�@��@�T= �c<��]>*��H>V>��3�>���J<���<�p�q�x���� �?� ��C�  <(�U��� 4Vr�33���@
���A@��? R�oD��mR�x���Q� �t����Z�Џ��؏��,��i?�7N�>��(�>�@Z�=�{��J��G�v�G�J�B�E�����a���@ǐ@���@~��@Q�?L *���ŲI�PP���&���'���@�K����Ag�q�PC��  C���C�uy�
���ʯ ?�7� ��?)6J��꡷ �
6t�V26tQ:6J�み)A D�Cj�ZD ��>(���4���X���v���*
�C3���5�2B���F�ǿB��ֿ�����E�t�.�����x= �W�����P����S�3ϔ�	CT�_CONFIG �K3����eg��STB_F_TTS��
����"�������{�M�AU���MSW�_CF��L  �K �OCVIEWf	�MI�U��� �߭߿��������� �0�B�T�f�x��� ������������,� >�P�b�t�������� ��������(:L ^p����� � �6HZl ~������,/��RCB�N��!�X.F/{/j/�/�/��/�/�/��SBL_�FAULT O�9*^�1GPMSK���7��TDIAG� P��U�����qUD1:� 6789012345q2�q���%P�ϭ?�?�?�?�?O O+O=OOOaOsO�O�O��O�O�O �a6�I'�
��?_��TRECPJ?\:
j4\_�7u[�? �_�_�_�_�_�_oo (o:oLo^opo�o�o�o��o�O�O_ _�UM�P_OPTION��>qTRB���9�;uPME��.Y�_TEMP  ?È�3B����ps�A�pytUNI'���ŏq6�YN_BR�K Qt�_�EDITOR q&qh�r�_2PENT 1R�9)  ,&�PEGA_BAR�RA_ESTEI�RA &p5� &�MAIN _P�LACE0 RV�IS$ra� &�PICK1Q����&COLOCA�_bpA_I�����&��PRENS�A ���&SGEGU(�%��P�p��  &-BCKEDT- (���pNO��o�PR�OG_1 /�A�SUMIR$�`�j��DROP_DEsFE�pX�ERT�������2������3��l���ANTEONA_C�m����SEM�� �o�Ф���o�E�x�UP��M������a�	�(ȯ*���F��DՆ���r��������p�
� �����J����pMG?DI_STA�u~���q�uNC_INF�O 1SI��b�������Կⷮ���;1TI� ��o#��|�G�d�o}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������Hu� �2�D� R�j�R�x������ ��������,�>�P� b�t������������� Z��#5Ga�k }������� 1CUgy� �������	// -/?/Yc/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?��?O%O7OQ/GO mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�?Oo o/o�_[Oeowo�o�o �o�o�o�o�o+ =Oas���� ��_�_��'�9�So ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�K�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�C� 5�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������ ���!�;�M�W�i�{� ������������� �/�A�S�e�w����� ����������+ E�Oas���� ���'9K ]o����1�� ��/#/=G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?��?�?	OO 5/?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�? �_�_oo-O#oIo[o moo�o�o�o�o�o�o �o!3EWi{ ����_�_��� �7oA�S�e�w����� ����я�����+� =�O�a�s�������� �ߟ���/�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������͟׿��� �'�1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ſ���������;� M�_�q������� ������%�7�I�[� m�������߯����� ���)�3EWi{ ������� /ASew�� �������/!+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?/��?�? �?�?/#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�?�_�_�_�_Oo -o?oQocouo�o�o�o �o�o�o�o); M_q���_�� ��	o�%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ����ß՟矝�� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߩ���������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u����߫� ����������); M_q����� ��%7I[ m�������� /!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�� �?�?�?�?�OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�?�?�_�_�_�_ �?�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy�_ �����_�	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q��y�����˟ �۟��%�7�I�[� m��������ǯٯ� ���!�3�E�W�i���� �$ENETM�ODE 1U���  
��������»���RROR_PRO/G %��%������TABLE  ���Q�c�u�����SEV_NU�M ��  �������_AU�TO_ENB  q̵��ݴ_NO��� V�������  *��������������+���(�<:���FLTR���ƇHIS�Ð�����_�ALM 1W��� ����̍�+ ;���������0�?߹_����  �����²u꒰TCP_�VER !��!���@�$EXTLO�G_REQv������SIZ����SkTK�������TOL  ��D�z~��A ��_BWDU�*�Z�V�ǲv?�DID� X敇Z�����[�S�TEPl�~�����O�P_DO���FA�CTORY_TU�Nv�d��DR_G�RP 1Y��`�d� 	p�.° ��*u���R�HB ��2 ���� �e9 ����bt� B�<�B�Q�C�P�Cj��BT�=C�]Ê�@��SA�Q��B2��A��A���BP[�� ����
C.�gR  A!~}�@��@.��u��
 JxO1�����-���o��_/�(/�	��  F!A�  @w�33R"�33�UUTn*@P  /�ȷ>u.�>*�߭<��ǊE��� F@ �"��5W�%�J��N�Jk�I'PK�Hu��IP�s�F!���?� � ?�/9�<9��896�C'6<,5�����Vv��7޷�t� ��� ��������FEATU�RE Z�V��ƱHand�lingTool� �5��Eng�lish Dictionary�7�4D St�0ar�d�6�5Analo�g I/O�7�7g�le Shift� Outo Sof�tware Up�date%Imat�ic Backu�p�9SAgroun?d Edit�0�7�Camera�0F��?CnrRndI�mXC�Lommon� calib U�I�C�FnqA�@Mo�nitor�Ktr~�0Reliab@��8DHCP�IZa�ta Acqui�s�CYiagno�sOA�1[ocum�ent View�e�BWual C�heck Saf�ety�A�6hanGced�F�:�UsnP�Fr�@�7xt. oDIO �@fiRT��Wend�PErr��@LQR�]�Ws�Yr��0�P E�:FCT�N Menu�Pv| S8gTP In'`�facNe�5Gig�E`nrej@p Ma�sk Exc�Pg��WHT^`Prox�y SvoT�fig�h-Spe�PSk�i�D�eJP�PmmuwnicN@ons�h�urE`'`_�1abc�onnect 2�xncr``str�u�2z>peeQPJ�QU�4KAREL �Cmd. L�`u�a�husRun-T�i�PEnvkx(`e�l +R@sP@S/�W�7Licens�e�Sn\�PBook�(System)��:MACROs,~�b/Offse@��uH�P8@_�pMR��@�BP^MechStop�at.p6R�ui�RKj�x�P�0P@�)�od@witc�h��>�EQ.���O�ptmЏ>��`fi�ln\=�gw�uul�ti-T�`tC�9P?CM funHwF��o3T�R?�f�Regei�pr�`I�rigP�FV����0Num �Selb����P Adju�`���J�tatu��
�iZ�5�RDM Robo}t�0scove�1�F�ea7��PFre�q Anly�gRem`��Qn�7F�R�Servo�P���8?SNPX b�rN;SN^`ClifQɮBLibr�3鯢0Q q�����o�ptE`�ssag?��4�� 0-C��;��/I_mB��MILIBk�E�P� Firm6BU�P�EcAcck@sKTPsTX_C�eln����F��1�V�orq}u@imula�A4�A�u��Pa�qU��j@�Ã&�`ev.�B�.@riP޿U�SB port ��@iP�PagP��R� EVNT�ϗ�n?except�P���t��ſX�]VC�Ar�b�bf�V2PҦ�$�4���SܠSCصV�gSGEk�a�UI�;?Web Pl!��ހ���Խ`�TeQfZDT Appl�d�:�ƺ� �GridV�play�R�WD
4�R
�.�:n�EQ+���r-10iA/7�L*��1Graph�ic���5dv�SD�CSJ�ck�q�5l�arm Caus�e/��ed�8As�cii�a��Loa9dnP�Upl,�Ol�0�AGu�6N�`���yFyc@�r������PV��Jo��m� �c�R���c���m�.�/�����Q�2*u:eR�AJ��P�ٶ4eqin8L����8NRT��9�On�0e Hel�HJ�`oI�alletiz?�H�����_��tr�[ROS E#th�q��T@e�ׅ��!�n�%�2D�tPk�g&Upg�~�(2DV-�3?D Tri-jQE�AưDef.qEBa)pdei��� �bImπF�f���nsp.q=�464MB DRAMZ�,#FRO5/@ell�<�Mshf!r/�'�c%3@pLƖ,ty@s˒xG��m��.[�� ��BU��8�Q�B�=mai�P߫В]Q����@q6wlu�����^`�xR�?eL� Sup������0�P�`cr��@�R����b䚮�pr1uest��rt~QQ��ߋL@!�4O��q$�K��_l Bui7�n��OAPLCOO�EVl%��CGU�OCRG��O��DR��O
TLSL_��BU/_��K�qLN_d�TA�OxVB�_��W�ܑZ���_TCB@�_�V�_�W���WF+o��V�O�W._�W�ņoTEH�o�f�O�gt�oTEj�xVF�_w�_xVGoTwBTw~oxVH�xVIA��v�&xVLN�yUMz��bo�f_xVN�xVP����^xVR&xVS��܇ʏ��W��v����VGF:�L�P2 _h��h�V�h��_g�	D��h�FFoh��g�sRD�� TUT���01:�L�2V�L�T�BGG��v�rai�n�UI��
%HM9I���pon��m�f�"�F�&�KAREL9� �T�Pj��<6 SWIoMESTڢF0O�<5�
"a�X�j����� ��ͿĿֿ���'�� 0�]�T�fϓϊϜ��� ��������#��,�Y� P�bߏ߆ߘ��߼��� ������(�U�L�^� ������������� ��$�Q�H�Z���~� ������������  MDV�z�� ����
I @Rv���� ��///E/</N/ {/r/�/�/�/�/�/�/ ???A?8?J?w?n? �?�?�?�?�?�?O�? O=O4OFOsOjO|O�O �O�O�O�O_�O_9_ 0_B_o_f_x_�_�_�_ �_�_�_�_o5o,o>o koboto�o�o�o�o�o �o�o1(:g^ p�������  �-�$�6�c�Z�l��� ������Ə����)�  �2�_�V�h������� ������%��.� [�R�d����������� ����!��*�W�N� `������������޿ ���&�S�J�\ω� �ϒϤ϶�������� �"�O�F�X߅�|ߎ� �߲���������� K�B�T��x���� ���������G�>� P�}�t����������� ��C:Ly p������	  ?6Hul~ �����/�/ ;/2/D/q/h/z/�/�/ �/�/�/?�/
?7?.? @?m?d?v?�?�?�?�? �?�?�?O3O*O<OiO `OrO�O�O�O�O�O�O �O_/_&_8_e_\_n_ �_�_�_�_�_�_�_�_ +o"o4oaoXojo|o�o �o�o�o�o�o�o' 0]Tfx��� ����#��,�Y� P�b�t���������� �����(�U�L�^� p����������ܟ� ��$�Q�H�Z�l�~� �������د���� �M�D�V�h��� � H552�}���21��R78���50��J614ީ�ATUPͶ54�5͸6��VCAMCRI�UIFvͷ28	�NRE���52��R63��S{CH��DOCV]�wCSU��869ͷ�0ضEIOC9�4R69��ESE�T���J7��R6�8��MASK��P�RXY!�7��OC�O��3帨���̸3��J6˸53��H�2�LCH��OPL�G�0�MHCR���S{�MCS�0���55ضMDSW����OP�MPR��M�@�0̶PCM �R0���ض��@�[51�51<�0�PRS��69�F{RD�FREQ���MCN��93̶S�NBAE�3�SHLEB��M��M���2̶�HTC�TMILܵ���TPA��TPTX��EL��Ѐ�q8������J95,ƷTUT�95�U�EV��UEC��U�FR�VCC��O��VIP�CSCN,�CSG8�r�I��wWEB�HTT䶳R6C�N�CGI�G��IPGS)R�C�DG�H77���6ضR85��R[66�R7��R:�R530�680�2��q�J��H�6<�6�,�RJح�0�4�6�o64\�5�NV�D��R6��R84�Tg����8�90l\���J93�91�b 7+���,�D0o�F�CLI���C�MS�� �STYF��TO�q���7ȻNN�ORS��J�% ��j�OL(EN�D��L��Sf(FV�R��V3D���P�BV,�APL��A�PV�CCG�C�CR|�CD��CD�L@CSBt�CS�K��CT�CTBL9��U0,(C��y0L8�C��TC �y0�'T�C(7TC��CTE\��07TEh��0���TFd8F,(GL8GI�8H�8I��E@�8�7�CTM,(M�8M�@8N�8PHHPL8R,d8(TSd8W�I@�VGF�GP2��P�2���@�H{7VPD��HF �VPSGVP�R�&VT��YP��VkTB7Vs�IH��VI aH'VK��VGene�����_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O?�a?s?�?  H55hT�1�1[Un�3R78�<50�9�J614�9ATU\�T�4545�<6�9�VCA�D�3CRIf,KUI8T�528-J�NRE�:52JR�63�;SCH�9D�OCV�JCU�48�69�;0�:EIOt�TsE4�:R69J�ESET�;KJ7�KR68�JMAS�K�9PRXYML7.�:OCO\3�<�J�)P�<3|ZJ6�<5u3�JH�\LCH\Z�OPLG�;0�ZM�HCR]ZSkMC�S�<0,[55�:MgDSW}k�[OP�[GMPR�Z�@�\0�:7PCMLJR0�k)P��:)`�[51K51�|0JPRS[6�9|ZFRD<JFR�EQ�:MCN�:9=3�:SNBA}K�[/SHLB�zM�{�@�ll2�:HTC�:T�MIL�<�JTPA��JTPTX�EL��z)`�K8�;�0�JJ�95\JTUT�[9�5|ZUEVZUE�C\ZUFR<JVCuC��O<jVIP,�wCSC\�CSGlJ��@I�9WEB�:H�TT�:R6{L��C�G{�IG[�IPGmS��RC,�DG�[�H77�<6�:R8�5�JR66JR7�[R|R53{6%8|2�Z�@Jml,|6|6\JR�\	P|�4L�6�64��5n�kNVDZR6+k�R84<���IP,�8f��90���KJ9�\91��̫7[KIP\J�D0�F��CLI�lKCMS�J9��:7STY,�TO�:�@��K7�LNN|ZOR�S<jJ��MZZ|OL�K�END�:L�S��FVR�JV3D�,�KKPBV\�AP�L�JAPV�ZCC�G�:CCRjCD��CDL̚CSBn�JCSK�jCTK��CTB��\���\�Ch�z���CL�TCLJl�l�TC��TCZ�CTE�J��|�TEX�J��<�TF��F\̥G��G��l�Hl�Ip�z)�l�k�CTM\�UM\�M��Nl�P,�eP��R��;�TS�ܹW��̚VGF��P2��P2�z ��VPDFLJVPn;�VPR��VT�;\� �JVTB��V�K�IH�VِM�<�V�K,�V{�Gene �8�83EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���� �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	- ?Qcu���� ���);M _q������ �//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�7}�0STD�4?LANG�4�9 �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2��D�V�RBT�6OPTNm��������Ǐ ُ����!�3�E�W��i�{�������ß�5DPN�4�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}ߏ�<�߳�ted �4�8 ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� �������������� );M_q�� �����% 7I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_o#o5o GoYoko}o�o�o�o�o �o�o�o1CU gy������ �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q����� ����˟ݟ���%� 7�I�[�m�������� ǯٯ������*��<�N�`�r���99����$FEAT_�ADD ?	��������  	��ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-?�Qcu�����D�EMO Z��   ���}� �'��0�]�T�f��� ������������#� �,�Y�P�b������� ����������(� U�L�^����������� �ܯ���$�Q�H� Z���~��������ؿ ��� �M�D�Vσ� zόϦϰ�������� 
��I�@�R��v߈� �߬���������� E�<�N�{�r���� ���������A�8� J�w�n����������� ����=4Fs j|����� �90Bofx �������/ 5/,/>/k/b/t/�/�/ �/�/�/�/�/?1?(? :?g?^?p?�?�?�?�? �?�?�? O-O$O6OcO ZOlO�O�O�O�O�O�O �O�O)_ _2___V_h_ �_�_�_�_�_�_�_�_ %oo.o[oRodo~o�o �o�o�o�o�o�o! *WN`z��� ������&�S� J�\�v���������� ڏ���"�O�F�X� r�|�������ߟ֟� ���K�B�T�n�x� ������ۯү��� �G�>�P�j�t����� ��׿ο����C� :�L�f�pϝϔϦ��� ����	� ��?�6�H� b�lߙߐߢ������� ����;�2�D�^�h� ������������� 
�7�.�@�Z�d����� ������������3 *<V`���� ����/&8 R\������ ���+/"/4/N/X/ �/|/�/�/�/�/�/�/ �/'??0?J?T?�?x? �?�?�?�?�?�?�?#O O,OFOPO}OtO�O�O �O�O�O�O�O__(_ B_L_y_p_�_�_�_�_ �_�_�_oo$o>oHo uolo~o�o�o�o�o�o �o :Dqh z������� 
��6�@�m�d�v��� ����ُЏ���� 2�<�i�`�r������� ՟̟ޟ���.�8� e�\�n�������ѯȯ گ����*�4�a�X� j�������ͿĿֿ� ���&�0�]�T�fϓ� �Ϝ������������ "�,�Y�P�bߏ߆ߘ� �߼���������(� U�L�^������� ������ ��$�Q�H� Z���~����������� ���� MDV� z������� I@Rv� ������// E/</N/{/r/�/�/�/ �/�/�/�/
??A?8? J?w?n?�?�?�?�?�? �?�?OO=O4OFOsO jO|O�O�O�O�O�O�O __9_0_B_o_f_x_ �_�_�_�_�_�_�_o 5o,o>okoboto�o�o �o�o�o�o�o1( :g^p���� ��� �-�$�6�c� Z�l�������ϏƏ؏ ���)� �2�_�V�h� ������˟ԟ��� %��.�[�R�d����� ��ǯ��Я���!�� *�W�N�`�������ÿ ��̿����&�S� J�\ωπϒϿ϶��� ������"�O�F�X� ��|ߎ߻߲������� ���K�B�T��x� ������������ �G�>�P�}�t�����|����  �� ����"4FXj |������� 0BTfx� ������// ,/>/P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�?�? �?�? OO$O6OHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t������� ��ο����(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz������y  �x�q���&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���� (�:�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p���(���q�p�x� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p��������������$FE�AT_DEMOIoN  �� ������INDE�X���IL�ECOMP [����B���8 SETUPo2 \BL?�  N w5�_AP2BCK �1]B	  �)����%����E �	���5� Y�f��B� �x/�1/C/�g/ ��/�/,/�/P/�/t/ �/?�/??�/c?u?? �?(?�?�?^?�?�?O )O�?MO�?qO O~O�O 6O�OZO�O_�O%_�O I_[_�O__�_�_D_ �_h_�_�_
o3o�_Wo �_{o�oo�o@o�o�o vo�o/A�oe�o ���N�r� ��=��a�s���� &���͏\�񏀏��� "�K�ڏo�������4� ɟX������#���G� Y��}����0���ׯtQ	� P� 2� *.VRޯ(���*+�Q���W�{�e���PC������F'R6:��ؾg�����T   �2����\�� ��d�*.F���ϕ�	ó����8o�ߓ�STM�9���ư%�d��ψߓ�HU߻�Jש�f�x����GIF�A�L�-�p���ߑ��JPG����Lձ�n�����JS�H�����6����%
JavaSc�riptt���CS�e���Kֹ�v� %�Cascadin�g Style ?Sheets��j��
ARGNAME�.DT'��O�\@;��[�k|(k DISP*rUO������ �
T�PEINS.XML/�:\Cc�Custom T?oolbar��	�PASSWORD����FRS:\��� %Pas�sword Config/c�Q/� J/�/���/:/�/�/p/ ?�/)?;?�/_?�/�? ?$?�?H?�?l?�?O �?7O�?[OmO�?�O O �O�OVO�OzO_�O�O E_�Oi_�Ob_�_._�_ R_�_�_�_o�_AoSo �_woo�o*o<o�o`o �o�o�o+�oO�os ��8��n� �'���]����� z���F�ۏj������ 5�ďY�k�������� B�T��x�����C� ҟg�������,���P� ��������?�ί� u����(���Ͽ^�� ���)ϸ�M�ܿqσ� ϧ�6���Z�l�ߐ� %ߴ��[����ߣ� ��D���h�����3� ��W����ߍ���@� ����v����/�A��� e������*���N��� r�����=��6s �&��\�� '�K�o� �4�X���#/ �G/Y/�}//�/�/ B/�/f/�/�/�/1?�/ U?�/N?�??�?>?�? �?t?	O�?-O?O�?cO��?�OO(O�O�F�$�FILE_DGB�CK 1]����@��� < �)
SU�MMARY.DG<�OsLMD:�O;_�@Diag Summary<_�IJ
CONSLO�G1__&Q_�_NQ�Console �log�_HK	TPOACCN�_o%o�?oJUTP Accountin�_�IJFR6:IP�KDMP.ZIP�sowH
�o�oKU[`E�xception��oyk'PMEMCH�ECK5o�_*_K��QMemory �DataL�F0�l�)6qRIPE�_$6�Zs%��q Packet� L�_�DL�$�<	r�qSTAT��|�S� %�r?StatusT��	FTP���:����Vw�Qmment� TBD؏� >�I)ETHERNE���
q�[�NQEthern�p~�Pfigura�o�ODDCSVRF�̏��ďݟd��� �verify asll��{D�.���DIFF՟��͟b�<�s��diffd��|
q��CHG01Y��@�R��f�z���-?��2ݯį֯k�v�����3a�H�Z��� ��ϥ�V�TRNDIAG.�LS�̿޿s�^q�3� Ope���q ~SQnosticEW���)VDEV7�DATt�Q�cϼu�g�Vis��D�evice�Ϫ�IMG7ºo����y��s=�Imagߨ�7UP��ES��T�?FRS:\�� ��OQUpdate?s List �IJ�g�FLEXEV�ENQ�X�j߃�f��F� UIF Ev����B,�s�)�
PSRBWLD'.CM��sL�������PPS_ROBOOWEL��GLo��GRAPHICS�4Dy�b�t��%�4D Grap�hics Filyeu��AOɿ�rGIG���u�
YvGigE�ة�B�N�? )��HADOW������\sShadow? Chang���v�bQRCME�RR�n�\s�� CFG Err{or�tail�� MA��CMSGLIB� �"^o� ��To�)�ZD��p��/XwZD6 �ad�HPNO�TI���
/�/ZuNotific��H/��AGUO�/yO ?�O'?P?OOt??�? �?9?�?]?�?O�?(O �?LO^O�?�OO�O5O �O�OkO _�O$_6_�O Z_�O~_�__�_C_�_ �_y_o�_2o�_?oho �_�oo�o�oQo�ouo 
�o@�odv �)�M���� �<�N��r������ 7�̏[������&��� J�ُW������3�ȟ ڟi�����"�4�ßX� �|������A�֯e� ����0���T�f��� �������O��s�� ϩ�>�Ϳb��oϘ� 'ϼ�K����ρ�ߥ� :�L���p��ϔߦ�5� ��Y���}���$��H� ��l�~���1����� g���� �2���V��� z�	�����?���c��� 
��.��Rd��� ��M�q� <�`���% �I��/�8/ J/�n/��/!/�/�/ W/�/{/?"?�/F?�/�j?|??�?/?�?�?��$FILE_FR�SPRT  ����0�����8MDONL�Y 1]�5�0� 
 �)MD�:_VDAEXTP.ZZZ�?�?_O�nK6%NO� Back fi�le 9O�4S�6Pe?�OOO�O�?�O_ _?>_�Ob_t__�_'_ �_�_]_�_�_o(o�_ Lo�_po�_}o�o5o�o Yo�o �o$�oHZ �o~��C�g ��	�2��V��z� �����?�ԏ�u�
��.�@��4VISB�CKHA&C*.�VDA�����FR�:\Z�ION\DOATA\v�����Vision VD�B��ŏ���'� 5��Y��j������ B�ׯ�x����1��� үg�������X���P� �t���Ϫ�?�οc� u�ϙ�(Ͻ�L�^��� ���)���M���q� � �ߧ�6���Z����߀%��I�������:L�UI_CONFIoG ^�5m�>�� $ h�F{�5������)�;�I���|xq�s����� ������a��� $ 6��Gl~��� K��� 2� Vhz���G� ��
//./�R/d/ v/�/�/�/C/�/�/�/ ??*?�/N?`?r?�? �?�???�?�?�?OO &O�?JO\OnO�O�O)O �O�O�O�O�O_�O4_ F_X_j_|_�_%_�_�_ �_�_�_o�_0oBoTo foxo�o!o�o�o�o�o �o�o,>Pbt ������� �(�:�L�^�p���� ����ʏ܏���$� 6�H�Z�l�������� Ɵ؟ꟁ�� �2�D� V�h���������¯ԯ �}�
��.�@�R�d� ����������п�y� ��*�<�N�`����� �ϨϺ�����u��� &�8�J���[߀ߒߤ� ����_������"�4� F���j�|������ [�������0�B��� f�x���������W��� ��,>��bt ����O���(:�  �xFS�$FLU�I_DATA �_������uRES�ULT 2`��� �T��/wizard/�guided/s�teps/Expertb��// +/=/O/a/s/�/�/�*��Contin�ue with =G�ance�/�/ �/??(?:?L?^?p?X�?�?�? T-U|��90 �� ��?���9��ps�?0OBOTOfOxO�O �O�O�O�O�O�O� � _/_A_S_e_w_�_�_ �_�_�_�_�_n�?�?t�?�<Frip� Oo�o�o�o�o�o�o �o!3E_i{ �������� �/�A�S�o$on�Ho�AO�Time?US/DST[�� ����+�=�O�a�s�������'Enabl�/˟ݟ���%��7�I�[�m������T�?{�ݯ����Æ24Ώ3�E�W�i�{� ������ÿտ翦��� �/�A�S�e�wωϛ� �Ͽ������ϴ�Ưد�� G��Region�χߙ߽߫��߀������)�;�+Americaso u�����������@��)�;��?�y��#߅�G�Y��ditorL�������#�5GYk}��+ �Touch Pa�nel �� (recommen�)���*<@N`r��U��e��w��������accesd�./@/R/d/v/��/�/�/�/�/�/Q|�Connect �to Network�/(?:?L?^?p? �?�?�?�?�?�?�?Y���������!�/��Introducts߆O�O�O�O �O�O�O__(_:_U ^_p_�_�_�_�_�_�_��_ oo$o6oHo  e�Oeo?O�X_�o�o �o�o'9K] o��R_���� ��#�5�G�Y�k�}�D����h`�ooj}o ߏ�o��*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ쯫��� Ϗ1��X�j�|����� ��Ŀֿ�����0� �A�f�xϊϜϮ��� ��������,�>��� _�!���E��߼����� ����(�:�L�^�p� ���߸������� � �$�6�H�Z�l�~��� O߱�s�������  2DVhz��� �����
.@ Rdv����� ���/��'/���`/ r/�/�/�/�/�/�/�/ ??&?8?�\?n?�? �?�?�?�?�?�?�?O "O4O�UO/yO�OO? �O�O�O�O�O__0_ B_T_f_x_�_I?�_�_ �_�_�_oo,o>oPo boto�oEO�OiO�o�o �O(:L^p �������_ � �$�6�H�Z�l�~��� ����Ə؏�o�o�o� /��oV�h�z������� ԟ���
��.�� R�d�v���������Я �����*����� ���C�����̿޿� ��&�8�J�\�nπ� ?��϶���������� "�4�F�X�j�|ߎ�M� _�q��ߕ�����0� B�T�f�x������ �������,�>�P� b�t������������� �߱���%��L^p �������  $��5Zl~� ������/ / 2/��S/w/9�/�/ �/�/�/�/
??.?@? R?d?v?�?�/�?�?�? �?�?OO*O<ONO`O rO�OC/�Og/�O�/�O __&_8_J_\_n_�_ �_�_�_�_�_�?�_o "o4oFoXojo|o�o�o �o�o�o�O�o�O�O �oTfx���� �����,��_P� b�t���������Ώ�� ���(��oI�m� �C�����ʟܟ� � �$�6�H�Z�l�~�=� ����Ưد���� � 2�D�V�h�z�9���]� ��ѿ����
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ��ߋ�տ ����#��J�\�n�� ������������� "���F�X�j�|����� ������������ ����u7��� ���,>P bt3������ �//(/:/L/^/p/ �/ASe�/��/ ? ?$?6?H?Z?l?~?�? �?�?�?��?�?O O 2ODOVOhOzO�O�O�O �O�O�/�/�/_�/@_ R_d_v_�_�_�_�_�_ �_�_oo�?)oNo`o ro�o�o�o�o�o�o�o &�OG	_k-_ �������� "�4�F�X�j�|���� ��ď֏�����0� B�T�f�x�7��[�� �����,�>�P� b�t���������ί�� ���(�:�L�^�p� ��������ʿ��뿭� �џӿH�Z�l�~ϐ� �ϴ���������� � ߯D�V�h�zߌߞ߰� ��������
��ۿ=� ��a�s�7ߚ����� ������*�<�N�`� r�1ߖ����������� &8J\n-� w�Q������ "4FXj|�� ������//0/ B/T/f/x/�/�/�/�/ ���/?�>?P? b?t?�?�?�?�?�?�? �?OO�:OLO^OpO �O�O�O�O�O�O�O _ _�/�/�/?i_+?�_ �_�_�_�_�_�_o o 2oDoVoho'O�o�o�o �o�o�o�o
.@ Rdv5_G_Y_�}_ ����*�<�N�`� r���������yoޏ�� ��&�8�J�\�n��� ������ȟ���� �4�F�X�j�|����� ��į֯����ˏ� B�T�f�x��������� ҿ�����ٟ;��� _�!��ϘϪϼ����� ����(�:�L�^�p� �ϔߦ߸������� � �$�6�H�Z�l�+ύ� Oϱ�s�������� � 2�D�V�h�z������� ��������
.@ Rdv����}� ������<N` r������� //��8/J/\/n/�/ �/�/�/�/�/�/�/? �1?�U?g?+/�?�? �?�?�?�?�?OO0O BOTOfO%/�O�O�O�O �O�O�O__,_>_P_ b_!?k?E?�_�_{?�_ �_oo(o:oLo^opo �o�o�o�owO�o�o  $6HZl~� ��s_�_�_���_ 2�D�V�h�z������� ԏ���
��o.�@� R�d�v���������П ��������]� ���������̯ޯ� ��&�8�J�\���� ������ȿڿ���� "�4�F�X�j�)�;�M� ��q���������0� B�T�f�xߊߜ߮�m� ��������,�>�P� b�t�����{ύ� �����(�:�L�^�p� ��������������  ��6HZl~� �������� /��S�z��� ����
//./@/ R/d/u�/�/�/�/�/ �/�/??*?<?N?`? �?C�?g�?�?�? OO&O8OJO\OnO�O �O�O�Ou/�O�O�O_ "_4_F_X_j_|_�_�_ �_q?�_�?�_�?�_0o BoTofoxo�o�o�o�o �o�o�o�O,>P bt������ ���_%��_I�[� ��������ʏ܏� � �$�6�H�Z�~��� ����Ɵ؟���� � 2�D�V��_�9����� o�ԯ���
��.�@� R�d�v�������k�п �����*�<�N�`� rτϖϨ�g������� ����&�8�J�\�n߀� �ߤ߶��������߽� "�4�F�X�j�|��� ��������������� ��Q��x��������� ������,>P �t������ �(:L^� /�A��e���� / /$/6/H/Z/l/~/�/ �/a�/�/�/�/? ? 2?D?V?h?z?�?�?�? o���?�O.O@O ROdOvO�O�O�O�O�O �O�O�/_*_<_N_`_ r_�_�_�_�_�_�_�_ o�?#o�?Go	Ono�o �o�o�o�o�o�o�o "4FXio|�� �������0� B�T�ou�7o��[o�� ҏ�����,�>�P� b�t�������iΟ�� ���(�:�L�^�p� ������e�ǯ��믭� ��$�6�H�Z�l�~��� ����ƿؿ����� � 2�D�V�h�zόϞϰ� �������Ϸ��ۯ=� O��v߈ߚ߬߾��� ������*�<�N�� r����������� ��&�8�J�	�S�-� w���c��������� "4FXj|�� _�����0 BTfx��[��� �����/,/>/P/ b/t/�/�/�/�/�/�/ �/�?(?:?L?^?p? �?�?�?�?�?�?�?� ���EO/lO~O�O �O�O�O�O�O�O_ _ 2_D_?h_z_�_�_�_ �_�_�_�_
oo.o@o RoO#O5O�oYO�o�o �o�o*<N` r��U_���� ��&�8�J�\�n��� ����couo�o鏫o� "�4�F�X�j�|����� ��ğ֟蟧���0� B�T�f�x��������� ү������ُ;��� b�t���������ο� ���(�:�L�]�p� �ϔϦϸ������� � �$�6�H��i�+��� O������������ � 2�D�V�h�z���]� ��������
��.�@� R�d�v�����Y߻�}� ���ߣ�*<N` r������� ��&8J\n� ��������/ ��1/C/j/|/�/�/ �/�/�/�/�/??0? B?f?x?�?�?�?�? �?�?�?OO,O>O� G/!/kO�OW/�O�O�O �O__(_:_L_^_p_ �_�_S?�_�_�_�_ o o$o6oHoZolo~o�o OO�OsO�o�o�O  2DVhz��� ����_
��.�@� R�d�v���������Џ ⏡o�o�o�o9��o`� r���������̟ޟ� ��&�8��\�n��� ������ȯگ���� "�4�F���)���M� ��Ŀֿ�����0� B�T�f�xϊ�I����� ��������,�>�P� b�t߆ߘ�W�i�{��� ����(�:�L�^�p� ������������ �$�6�H�Z�l�~��� �������������� /��Vhz��� ����
.@ Qdv����� ��//*/</��]/ �/C�/�/�/�/�/ ??&?8?J?\?n?�? �?Q�?�?�?�?�?O "O4OFOXOjO|O�OM/ �Oq/�O�/�O__0_ B_T_f_x_�_�_�_�_ �_�_�?oo,o>oPo boto�o�o�o�o�o�o �O�O%7�_^p ������� � �$�6��_Z�l�~��� ����Ə؏���� � 2��o;_���K�� ԟ���
��.�@� R�d�v���G�����Я �����*�<�N�`� r���C���g���ۿ�� ��&�8�J�\�nπ� �Ϥ϶����ϙ���� "�4�F�X�j�|ߎߠ� �����ߕ�����˿-� �T�f�x������ ��������,���P� b�t������������� ��(:���� A�����  $6HZl~=� ������/ / 2/D/V/h/z/�/K] o�/��/
??.?@? R?d?v?�?�?�?�?�? ��?OO*O<ONO`O rO�O�O�O�O�O�O�/ �O�/#_�/J_\_n_�_ �_�_�_�_�_�_�_o "o4oE_Xojo|o�o�o �o�o�o�o�o0 �OQ_u7_��� �����,�>�P� b�t���Eo����Ώ�� ���(�:�L�^�p� ��A��eǟ��� � �$�6�H�Z�l�~��� ����Ưد����� � 2�D�V�h�z������� ¿Կ�������+�� R�d�vψϚϬϾ��� ������*��N�`� r߄ߖߨߺ������� ��&��/�	�S�}� ?Ϥ����������� "�4�F�X�j�|�;ߠ� ����������0 BTfx7��[� ����,>P bt������� �//(/:/L/^/p/ �/�/�/�/�/��� �!?�H?Z?l?~?�? �?�?�?�?�?�?O O �DOVOhOzO�O�O�O �O�O�O�O
__._�/ �/?s_5?�_�_�_�_ �_�_oo*o<oNo`o ro1O�o�o�o�o�o�o &8J\n� ?_Q_c_��_��� "�4�F�X�j�|����� ��ď�oՏ����0� B�T�f�x��������� ҟ����>�P� b�t���������ί� ���(�9�L�^�p� ��������ʿܿ� � �$��E��i�+��� �ϴ���������� � 2�D�V�h�z�9��߰� ��������
��.�@� R�d�v�5ϗ�Yϻ�}� �����*�<�N�`� r��������������� &8J\n� ��������� ��FXj|�� �����//�� B/T/f/x/�/�/�/�/ �/�/�/??�#� G?q?3�?�?�?�?�? �?OO(O:OLO^OpO //�O�O�O�O�O�O _ _$_6_H_Z_l_+?u? O?�_�_�?�_�_o o 2oDoVohozo�o�o�o �o�O�o�o
.@ Rdv����}_ �_�_�_��_<�N�`� r���������̏ޏ�� ���o8�J�\�n��� ������ȟڟ���� "����g�)����� ��į֯�����0� B�T�f�%��������� ҿ�����,�>�P� b�t�3�E�W���{��� ����(�:�L�^�p� �ߔߦ߸�w����� � �$�6�H�Z�l�~�� ������������ 2�D�V�h�z������� ��������
-�@ Rdv����� ����9��] �������� //&/8/J/\/n/- �/�/�/�/�/�/�/? "?4?F?X?j?)�?M �?qs?�?�?OO0O BOTOfOxO�O�O�O�O /�O�O__,_>_P_ b_t_�_�_�_�_{?�_ �?oo�O:oLo^opo �o�o�o�o�o�o�o  �O6HZl~� ��������_ o�_;�e�'o������ ԏ���
��.�@� R�d�#��������П �����*�<�N�`� �i�C�����y�ޯ� ��&�8�J�\�n��� ������u�ڿ���� "�4�F�X�j�|ώϠ� ��q�������	�˯0� B�T�f�xߊߜ߮��� �������ǿ,�>�P� b�t��������� ����������[�� ��������������  $6HZ�~� ������  2DVh'�9�K�� o����
//./@/ R/d/v/�/�/�/k�/ �/�/??*?<?N?`? r?�?�?�?�?y�?� �?�&O8OJO\OnO�O �O�O�O�O�O�O�O_ !O4_F_X_j_|_�_�_ �_�_�_�_�_o�?-o �?QoOxo�o�o�o�o �o�o�o,>P b!_������ ���(�:�L�^�o �Ao��eog�܏� � �$�6�H�Z�l�~��� ����s؟���� � 2�D�V�h�z������� o�ѯ�����˟.�@� R�d�v���������п ����ş*�<�N�`� rτϖϨϺ������� �����/�Y���� �ߤ߶���������� "�4�F�X��|��� ������������0� B�T��]�7߁���m� ������,>P bt���i��� �(:L^p ���e�w������ ��$/6/H/Z/l/~/�/ �/�/�/�/�/�/� ? 2?D?V?h?z?�?�?�? �?�?�?�?
O��� OO/vO�O�O�O�O�O �O�O__*_<_N_? r_�_�_�_�_�_�_�_ oo&o8oJo\oO-O ?O�ocO�o�o�o�o "4FXj|�� __������0� B�T�f�x�������mo Ϗ�o�o�,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � ��!��E��l�~��� ����ƿؿ���� � 2�D�V��zόϞϰ� ��������
��.�@� R��s�5���Y�[��� ������*�<�N�`� r����g������� ��&�8�J�\�n��� ����c����������� "4FXj|�� �������0 BTfx���� ���������#/M/ t/�/�/�/�/�/�/ �/??(?:?L?p? �?�?�?�?�?�?�? O O$O6OHO/Q/+/uO �Oa/�O�O�O�O_ _ 2_D_V_h_z_�_�_]? �_�_�_�_
oo.o@o Rodovo�o�oYOkO}O �O�o�O*<N` r������� �_�&�8�J�\�n��� ������ȏڏ����o �o�oC�j�|����� ��ğ֟�����0� B��f�x��������� ү�����,�>�P���!�3������$F�MR2_GRP �1a���� �C4  �B�[�	 [��߿�ܰE�� Fw@ 5W��S�ܰJ��NJk��I'PKHu���IP�sF!{���?�  W��S�ܰ9�<9��896C�'6<,5�{��A�  ��6��BHٳB�հ��޷�@�33�3�3S�۴��ܰ@UUT'�@��8���W�>u.�>*�߭<����=[��B=���=�|	<�K�<��q�=�mo����8�x	7H�<8�^6�?Hc7��x?��� �������"��F�X����_CFG b»T Q���|��X�NO º/
F0�� ��W��RM_CHKTYP  ��[�ʰ̰܂���ROM�_MsIN�[���9�u���X��SSBh��c�� ݶf�[�]����^��TP_DEF_O��[�ʳ��IR�COM���$G�ENOVRD_D�O.�d���THR�.� dd��_E�NB�� ��RA�VC��dO�Z�� ���Fs  G�!� GɃ�I��C�I(i J����+���%������ �QOUU��j¼������<6�i�C��;]�[�C� � D�+��@���B����.��R SMT��k�_	ΰ\��$HO7STCh�1l¹[���d�۰ MC�[���/Z��  27.0� 1�/  e�/?? '?9?G:�/j?|?�?�?��,Z?T3	anonymouy �?�?	O@O-O?N�/ڰRHRK �/�?�O�/�O�O�O�O _V?3_E_W_i_�O&_ �?�_�_�_�_�_@O�_ dOvOSo�_�Ojo�o�o �o�o_�o+= `o�_�_����� o&o8oJoL9��o]� o��������oɏۏ� ���4�j+�Y�k�}� �������� �� T�1�C�U�g������� ����ӯ��x�>��-� ?�Q�c�����Ο��� Ͽ����)�;ς� _�qσϕϧ�ʿ �� ����%�7�~����� ߶ϣ���������� �Ϻ�3�E�W�i�ߍ� �ϱ���������@�R� d�v�x�J��߉����� �������+= `���������:$h!ENT 1m� P!V  7 ?.c &�J�n��� /�)/�M//q/4/ �/X/j/�/�/�/�/? �/7?�/?m?0?�?T? �?x?�?�?�?O�?3O �?WOO{O>O�ObO�O �O�O�O�O_�OA__ e_(_:_�_^_�_�_�_��ZQUICC0 �_�_�_?od1@oo.o�od2�olo~o�o�!ROUTER��o�o�o/!PC�JOG0!�192.168.�0.10	o�SCA�MPRT�\!bpu1yp��vRT�o���� !So�ftware O�perator Panel�mn���NAME !~�
!ROBO��v�S_CFG 1�l�	 ��Auto-st�arted'�FTP2��I�K2� �V�h�z������� ԟ����	���@�R� d�v���	������ �:���)�;�M�_�&� ��������˿�p�� �%�7�I�[��"�4� F�ڿ��������!� 3���W�i�{ߍߟ��� D���������/�v� �Ϛ�w�ߛ��Ͽ��� ������+�=�O�a� ��������������� 8�J�\�n�p�]�� �������� #5X�k}�� ��0/D1/ xU/g/y/�/RH/�/ �/�/�//?�/??Q? c?u?�?���/? �?:/O)O;OMO_O&? �O�O�O�O�O�?pO_ _%_7_I_[_�?�?�? t_�O�_O�_�_o!o 3o�OWoio{o�o�_�o Do�o�o�o����_ERR n���-=vPDUSIZW  �`^�P�Tt�>muWRD ?�΅�Q�  guest�f�������~�S�CDMNGRP �2o΅WpC��Q�`���fKL�� 	P01.0�5 8�Q   ��|��  };|��  z[� ���w����*���Ť�x����[ݏȏ�V�בPԠ���~���)����D�Yr���؊p"�P�l�P���Dx��d�x�*�����%�_GR�OU7�pLyN���	/�o���QUP���UTu� �T�YàL}?pTT�P_AUTH 1�qL{ <!i?Pendan�����o֢!KAR�EL:*�������KC��ɯۯ��V�ISION SET�9����P�>�h� �f����������ҿ�����X�CTRL rL}O�uſa�
��mFFF�9E3-ϝTFR�S:DEFAUL�T��FANU�C Web Server�ʅ�t�X� ��t@���1�C�U��g�;tWR_CON�FIG s;� ���=qIDL_�CPU_PC���aBȠP�� BH���MIN�܅q��GNR_IOFq{r�`�Rx��NPT_SI�M_DO��S�TAL_SCRN�� �.�INTPMODNTOLQ����RTY0����-�\�ENBQ�-����OLNK 1tL{�p������)��;�M���MASTE��%���SLAVE� uL|�RAM�CACHEk�c�O>^�O_CFG�������UOC�����CMT_OP���Pz�YCL������_A�SG 1v;��q
 O�r���� ���&8J�\W�ENUMzs�Py
��IP����R?TRY_CN��PM�=�zs���Tu ������w���p/�p���P_MEMBE�RS 2x;�l� 5$��X"��?�Q'�W/i)��RCA_A�CC 2y� � X�P� ��� �  /�� 6��a&�� ��&4� �p�/�$  s��`�,�$�BUF001 2�z�= L�u0  u0L�:4��:4�:3M	R4�R4)R49R4JR4Z�R4kR4{R4�R4��R4�R4�u0p�]�M�u048�@�N:3N+u�0@5(NBu�0-0H Nbu�0:1N��4�u0�B�2�N��4�Z�4�:3ODD�&D6DHD�4O�m:3P g�@�YXP"u0^hg�Py0:1PqRD��u0)�K�P{�4u�48c�:3sc�rD�4K�e���e�K��D��D���DЂD�D�:4�:4:4#:42:4C*:4S:4d:4s:4�02<2�:4�4L�:392$?63:1@1ERI0ER Q0:1X1]Ra0]Ri0]R q0]RQD�1]R�0]R�0�]R�0d8��1g�8�1]R�0]R�0�A�3��1t� =`�1`�X�1�2��?0B03 �9Nx&� A:1Ab@ b@b!@b)@b�Tx8ATBA@g �HA TBQOSCi@jApA:1xAx}b�T�Ad� ؐA�Z���As�8�A�b�@�b�@�b�@ ER�@ER�@ER�@ER�@ ER�@ER�@ER�@ER�@ ER�4QER�0ERP:193-_65GSNrI2WS ��X3gSfri2wSfry2 �Sfr�2�Sfr�2_P�2 _P�2�Sfr�0���3�0 �0�r�0�r�P�rR�3 �r�2�0�2�0Bc� Bc�!B/c��t8C GcN�I@N��tXAN�a@ N�iBwc~�yB�c���C �`�B�`�B�`�B�c�� �B�cNr�B�cNr�B�c Nr�B�cNr�B�cNr�t�SsNrR6��2{��4r�}ŋ���<�����o�o��2�HIuS!2}� ܷ!� 2024-0'7-2�����Пp���GaQ�7 � N���*�<�N�`�o�X�cȩ�O���p����ɯ �  ;� ��`��" *c� N��"��,�>�.u��b꩘2��~������������m�b��l�����r��f=n��6-27m�Z�`l�~�ٯ��fnۿ����������"�g=�6I�6�H�Zߑ�o��o���g�Ϥ߶�8�����"�j�=ȴ�P�#�5������h��j��|���\��y��cN=�1���������� 9 ��cNw�\�n��� ����,P������������9� _� 1 Oas�s������(���,r�J�N�Qc����:� d� ;M_M�_����(��˶;3�bٰo� )/(/:/q:ϕ�/��/�/ �dd ��/�/ ??$?�$� Z?l?~?���"��"�% ���/�?�?�? O���� 6OHOZO�/�#:��% m��"u��"hO�O�O�O �����O_1_C_U��B�B a�%I�O�_ �_�_�_��5p����_o$o6o��!n���_o qo�o�o�o�O�o�o� ��b0t� ��AsN`r�r�@�o����˶�q ٰ�*�<�N�`�N/`/ �����̏���0� ���&��%�7�I�7? I?�����ڏ쏐�� ���%�O�_[�m��$�3t�����m� �u�ޟӯ����O�O R�?�Q�c�,�3t~�
�CrN���������п�_�RI_CFG� 2~�[ H�
Cycle T�ime(�Bu�sy�Idl��-�mi����S�Up� ��Read(�DCowG�C�bPX���Count �	N'um �.������(�����PROG����U�P��)/softpa�rt/genli�nk?curre�nt=menup�age,1133,1�C�U�g�y�T����SDT_ISO�LC  �Y� ����J23_D�SP_ENB  ���2���INC ����(���A  � ?�  =�̟�<#�
���:�o �2�D�(�X/�l���OB��C���O��ֆ�G_GR�OUP 1���}�2< ���P����t�?����(�Q'�L�^�p�/� ���������\�~��G_IN_AUT�O����POSRE����KANJI_�MASK0��DR�ELMON ��[��(�y���������f�Ã�����(�-��KCwL_L NUM���G$KEYLOGOGINGD�P�rQ�����LANGUA_GE �U���DEFAUgLT ��QLG������S��(�x��  8T�H�  �(�'0縤�(��Aߍ�;���
*!(UT1:\ J/ L/Y/k/ }/�/�/�/�/�/�/�/�$>(�H?�VLN_DISP ����P�&�$�^4OCTOL��Dz����
�1�GBOOK ���uQ1V�11uP ^P*O!O3OEOWOiK`yM�TËIgF	�5�)����O}���2_BUFF 2���G ~�[�u_ tR��6_M�R_d_�_�_ �_�_�_�_�_�_o3o *o<oNo`o�o�o�o�o����ADCS � �����L�O��+�=Oa�dIO 2��k ����������� ��*�:�L�^�r��� ������ʏ܏����$�6�J�uuER_ITM��d������ǟ ٟ����!�3�E�W� i�{�������ïկ�p����7x�SEVD���t�TYP�����s������)RS�Te�eSCRN__FL 2��}�����/�A�S�eόwϨ�TP{��b�>�=NGNAM��Eܮ�dUPSf0GI���2����_L�OAD��G %���%DROP_~�EITO_3�����MAXUALR�Mb2�@���
�K���_PR��2  h�3�AK�Ci0���qO=_'X�Ӭ�P 2]��; �*V	��-��
*����4 ��*��'�`�	xN�� z����������� 1�C�&�g�R���n��� ��������	��? *cFX���� ���;0 q\������ �/�/I/4/m/X/ �/�/�/�/�/�/�/�/ !??E?0?i?{?^?�? �?�?�?�?�?�?OO�AOSO6OwObO�OD�D;BG*� ��գ���ѤO�@_LDXD�ISA����ssME�MO_AP��E {?��
 �A x$_6_H_Z_l_~_�_��_K�FRQ_CF�G ����CAM w@��S�@<�ԃd%�\o�_�P�Ґ�����*Z`/\b **: eb�DXojho�F�o�o �o�o�o�o;�O ��dZ�U�y|��z,(9�Mt��� 1��B�g�N���r��� �����̏	���?�~A�ISC 1���K` ��O�����O����O֟����K�]�_M?STR �3���SCD 1�]� �l��{�����د ïկ���2��V�A� z�e�������Կ���� ���@�+�=�v�a� �υϾϩ�������� �<�'�`�K߄�oߨ� �ߥ��������&�� J�5�Z��k����� ����������F�1� j�U���y��������� ����0T?x6�MK�Q�,��Q��$MLTARM��R�?g� �~s�@���@ME�TPU�@l���4�NDSP_AD�COL�@!CM3NT7(FNSW�iSTLIx *%� �,�����Q��*POSC�F��PRPMlV�ST51�,�w 4�R#�
g! |qg%w/�'c/�/�/�/ �/�/�/?�/?G?)? ;?}?_?q?�?�?�?�?��1*SING_C�HK  {$M7ODA�S�e����#EDEV 	��J	MC:WLHOSIZE�Ml �#ETASK %�J�%$123456�789 �O�E!GT�RIG 1�,� l�Eo#_�y_S_��}�FYP�A�u9D�"CEM_INF �1�?k`)�AT&FV0E0�X_�])�QE0V�1&A3&B1&�D2&S0&C1�S0=�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_ �_o�3o��o�� �o��"�4��X� ��ASe֏�� �C�0���f�!��� q�����s�䟗����� ͏>��b���s���K� ��w���ٯ�ɟ۟ L����#�����Y�ʿ ����$�߿H�/� l�~�1���U�g�y��� �ϯ� �2�i�V�	�z��5ߋ߰ߗ���PONIwTOR�G ?kK�   	EX�EC1o�2�3��4�5��@�7*�8�9o�� ����(��4��@� ��L��X��d��p⨂�|��2��2��2���2��2��2��2���2��2��2��3ʉ�3��3(�#AR_�GRP_SV 1ݛ�[ (�1?������{b?�7N��b�?�=.IRM�A�_DsҔN��ION�_DB-@�1Ml/  �# �FH"�� �/� � �FH��N  � %�@%d�2��� �JE-ud1�}E���)PL_NAME !�E�� �!Def�ault Per�sonality� (from FsD)b (RR2��� 1�L�XL��p�X  d�-?Qcu� ������// )/;/M/_/q/�/�/�/EC2)�/�/�/??@,?>?P?b?t?EB<�/ �?�?�?�?�?�?
OO�.O@OROdO��6D�?�N
�O�O�P�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ �O�O2oDoVohozo�o �o�o�o�o�o�o
 .@o!ov��� ������*�<��N�`�r����� �Fs  GT��G�M���  #�ÏՍ�d���� ���(�6������
� �m�~�h����� ������ğ֟������:���
�]�m����	`������į��:�oA������ A�  /���P����r��� ����^�˿ݿȿ��t%��R�� 1��	�X ��, �� ��� a� @D7�  t�?�z�`��?� |��A/��xt�+��;�	l���	 �x7J���� � ^�� �<�@����� ��·�K���K ��K=*��J���J���J9��
��ԏC߷�@�t�@w{S�\��(Eh�����.��I����ڌ���T;�f�ґ�$��3���´  �@��>��Թ�$�  >�����ӧU���3x`���� �
�����Ǌ��� ��  {  @�T�����  ��H R n�ϊ�-�	'�� � ��I�� �  ��<�+�:�È����=�����0Ӂ���N �[��n @���f���f��k���,�av�  �'��Yэ�@2�?�@�0@�Ш����C��Cb C�G�\C������G��@�� �I ����� )�B�b $/�!��L�Dz�o�ߓ~���0��( �� -���������!9�D�  �9�恀?�ff0G�*<� }�qD�1�89��>��Hbp��(�(9��P���	������>�?�՚9�x9�W�<
�6b<߈;����<�ê<�?��<�^��I/2��A�{��fÌ¾,�?fff?_�?y&� T�@�.�"�J<?�\��"N\�5���!��(� |��/z��/j'��[0? ?T???x?c?�?�?�?`�?�?�?5��%F� �?2O�?VO�/wO�)IO��OEHG@ G@�09�G�� G} ଙO�O�O_	_B_-_\f_Q_BL9�B��Aw_[_�_b��_�[�_ ��mO3o�OZo�_~o�ox�o�o���b��PV( @|po	lo- *cU�ߡA���r59�CP�Lo�}?����#���5��W9���6�Cv�q�CH3� j�t�����q�����|^(�hA� �AL�ffA]��?��$�?��;����u�æ�)��	ff��C��#�
���g\)��"�33C�
������<��؎G�B����L�B�s?����	";��H�ۚG��!�G��WIY�E���C�+��8�I۪I�5��HgMG��3E��RC�j�=x�
�pI����G��fIV=�E<YD�C <�ݟȟ����7�"� [�F��j�������ٯ į���!��E�0�i� T�f�����ÿ���ҿ ����A�,�e�Pω� tϭϘ��ϼ������ +��O�:�s�^߃ߩ� ���߸������ �9� $�6�o�Z��~��� ���������5� �Y� D�}�h�����������@����
C.(�g���/"���<��t��q�3�8����q4�Mgu���q�V�wQ�
4p�+4�]$$dR��v���uPD"P��Q�_/Z/=/(/a/L+Rg/n/�/��/�/�/�/  %� �/�/+??O?:?s?/`�_�?�?�?�;�?��?O�? OFO4O�r LO^O�O�O�O�O�O�J  2 Fs�w�GT�V�MuBO�|r�pp�C��S@�R_�poy_�_؝_�_o \!�WɃh_oo(o�z�?���@@�zJ�D�p�pk1�p�~
 6o�o�o �o�o�o�o);�M_q�ڊsa �����D��$�MR_CABLE� 2�� )]��T�LaMaa?�PMaLb�p�Z�ɴ&P�C�p?aO4�>�B���?b��>?`F�ڈ�F�?b��v�_l  ��&P�v�^wdN�{0�_��V��R3���F�[�7�I�X�T��6P?`C$��Č���y�2�?`j&����F.S�,���| ��&Pr��C���=�����$��?`Z�RK�{F�h څ��s9�"T�p�� J�D�V�h�z�ߟڟ�� ��ԟ�K�
��F�@��R�d��	j��#?` ��������?b���A_N�`�r��?b*��** ��sOM ��y����{e`� ���%% 2345678901ɿB۵ ƿ���?`�?`j=�?`?a
��z�not segnt ���W��TESTFE�CSALG� egD�Z=�d��ga%�
���@��?d�r���������� 9U�D1:\main�tenancesG.xmS�.�@�vj��DEFAU�LT�\�rGRP {2���  p�R��I?e  �%1�st mecha�nical chgeck�?a���#������E��Z��(�:�L�^�?b��c�ontrolleAr�Ԍ��߰��D������ ��$�s�M��L�?b"8b���v��B�����������/�C}�a�6����dv���s��C��ge��. b?attery�&��E	S(:L^�p�	|�duiz�awblet  D�� ��љѿ�E���/"/4/s��g�reas�>gf�Br#-?`|!�/�E�@�/�/�/�/�/s�
��oi,�g/y/�/��/t?�?�?�?�?s�H�
�?f�W��1<?`AO�E
c?8OJO\OnO�O�t��?O��'O�O_ _2_D_s��OverhaulE��L��R x?`�Q�_���O�_�_�_�_o?`$�_0oϤFi 4oVٰ_�o�o�o�o�o o�o@oRodo%K] o���o�* ��#�5�G��X�}� ����ŏ׏���� \�1�C���g������� ����ӟ"���F�X�-� |�Q�c�u�����蟽� ���B��)�;�M� _�����ү䯹��ݿ ���%�t�IϘ��� �ο�ϵ�������:� �^�pςϔ�i�{ߍ� �߱� ���$�6�H�	� /�A�S�e�w��ߛ��� ���������+�z� <�a���d�������� ����@�'v�K�� o�����* <`5GYk} ����&�/ /1/C/�g/���/ ��/�/�/�/	?X/-? |/�/c?�/�?�?�?�? �??�?B?T?f?x?MO _OqO�O�O�?�OOO ,O�O_%_7_I_[_�O _�O�O�O�_�_�_�_8o!o�T	 T"oOo aoso�_�o�_�k�o�o �o�o�o�o2D z��`r��� ��.�@���v��� ��\�n�Џ⏤�����R ��Q?� ; @eQ �oW� i�{�eVC�����̟aXw*�**  � ����� �2�D��h�8z��������_�S ������կ7�I� [�����ɯ/���ǿٿ #���!�3�}����� {ύϟ��s������� C�U�g��S�e�w�9�@�߭߿�	��eUeQ��$MR_HIS�T 2������ 
 \jR$ 2�34567890�1*�2����)�9 c_���R��a_���� �����=�O�a��*� x�����r����� ��9��]o&�J �����#� G�k}4�Z��SKCFMAP � �������Z��ONREL  �����лEXC/FENB'
���!FNC$/$JO�GOVLIM'd��m �KEY'zp%y%_PAN(��"�"�RUN`,�p%�SFSPD�TYPD(%�SI�GN/$T1MO�Tb/!�_CE_GRP 1����"�:`��n?Z [?�?�؆?�?~?�?�? �?!O�?EO�?:O{O2O �O�OhO�O�O�O_�O /_�O(_e__�_�_�_ �_v_�_�_�_o�׻QZ_EDIT4���#TCOM_C_FG 1��'%�to�o�o 
Ua_A�RC_!"��O)T�_MN_MODE�6�Lj_SPL��o2&UAP_CP�L�o3$NOCHE�CK ?� � Rdv� ���������*�<�N�`��NO_?WAIT_L 7Jg650NT]a���UzZ��_ERR?12���ф��	���-����R�d����`O�����| ���
aB����o����C���������,V<� �� ?��Uϟj����قPA�RAMႳ��N�oR�=��o��� = e������ گ�ȯ��"�4��X�j�F�<�蜿��A��ҿ�"ODRDSP��c6/(OFFSET_CAR@`�o��DIS��S_A��`ARK7KiOPEN_FILE4��1�aKf�`OPTION_IO�/�!���M_PRG %��%$*����h�WmOT��E7O�����Z��  ���"�÷"�	� �V"�Z����RG_DSBOL  ��ˊ����RIENTT5O ZC����A �U�`IM_ED���O��V�?LCT ���Gb�ԛa�Zd��_P�EX�`7�*�RAT��g d/%*��UOP ���{��������������$�PAL�������_?POS_CHU�7�����2>3�L��XL�p��$�ÿU�g�y����� ����������	- ?Qcu����Y2C���"4 FXj|��� ��� //$/6/H/ Z/l/~/�Y���.��/�/ςP�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO�/�/ LO^OpO�O�O�O�O�O �O�O __$_6_H_Z_ )O;O�_�_�_�_�_�_ �_o o2oDoVohozo`�o�o�_<���o �m ���(�"{B Pw�m�m���~�jw8��w����� �2�T��p��w���H��t	`���̏ޏ��:�o����� �|2��pA�  I� �j�`�������� �џ���@��#��)�Or�1��_�� 8���, �\Ԡ��� @D�  ��?����~�?� ���!D�������%G�  �;�	l��	 ��xJ�젌����� ��<� ��� ���2�H(��H3�k7HSM5G��22G���GN�3%�R��oR�d�2�KCf��a��{�ׄ������/��3������4��>���К������3�A�q���{q�!ª��ֱ� "�(«�=ø2����� ��{�  @�Њ���/  ��Њ�2����.�	'� �� ��I� ��  �V�,�=�������˖ß����  �y��n @"��]�<߼+�������-�N�Д� C '�Ь�w�ӰC��C��\C߰������ߤ!���@��4���/��2�~�B���B�I�;�)�j客z +���쿱����������( �� -��#�����L��!�]�9�� > q�?�ffaH�Z��� ��������8� ����>�|P��}�(� ��P�����x��\�?��� �x� ���<
6b�<߈;܍��<�ê<����<�^�*�gv�A�)ۙ�脣��F�?offf?}�?&� ���@�.��J�<?�\��N\��)�������� ���ޤy�N9r ]������� /&/�J/5/n/��	g/�/c(G@ �G@0i�G�� G}���/??<?'?p`?K?�?o?BLi�B��A�?y?�?|��? K�?ů�/QO�/xO�?��O�O�O�Om��b�9�n�t @|�O'_��OK_6_H_�_lS��A��RS�i�Cn_�_j_<0O�]?��oo�Ao,o¹�Wi���fToC���`CHQo�>Jd�`a�a@I�ܚ>(hA�� �ALffA]���?�$�?����ź°u�����)�	ff��C�#�
�o�pg\)��33�C�
������<��nG��B���L��B�s�����	0źH�ۚ�G��!G��W�IYE����C�+�½I���I�5�Hg�MG�3E���RC�j=�~
��pI���G���fIV=�E<YD�#Zo��� 
��U�@�y�d����� ����я�����?� *�c�N���r������� �̟��)��9�_� J���n�����˯��� گ�%��I�4�m�X� ��|���ǿ���ֿ� ��3��W�B�Tύ�x� �Ϝ���������	�/� �S�>�w�bߛ߆߿� �߼�������=�(�ta�L�(q���)����Z�������a3�8�x�����a4Mgu��<���a�VwQ�(��4p�+4�] B�B���p���������J�UPbP���QO�%x�1[FjR�������  C���I4 mX�8
O������.//>/d/R/�Rj/|/�/�/��/�/�/:  2 �Fs�gGT�.&6�M�eBmp�R,�P�aC��3@�_p?��?�?�?�?�?�=�S��OO)O;OMO�c?_���@@�j���`�`�1�`�^
 TO�O�O�O �O�O_#_5_G_Y_k_�}_�_�_�j�A �����D��$P�ARAM_MEN�U ?B���  �DEFPULSE�{	WAITT�MOUTkRC�Vo SHE�LL_WRK.$�CUR_STYLv`DlOPTZ1NZoPTBooibC?oR_DECSN` ���l�o�o�o &OJ\n�������QSSREL?_ID  >�
1���uUSE_PR_OG %�Z%�@��sCCR` �
1��SS�_HOST !�Z!X���M�AT _���x�����|�L�_TIMEb� �h��PGDEB�UG�p�[�sGINP_FLMSK��E�T� V�G�PGA�r� 5��?��CH�S�D�TYPE�\�0��
�3�.�@� R�{�v�����ï��Я ����*�S�N�`� r����������޿� �+�&�8�J�s�nπ���ϻ�G�WORD �?	�[
 	�PR2��MAI��`�SU�a��T1EԀ���	Sd҇COL��C߸�LV� C�~�h��d*�TRACEC�TL 1�B���Q �� �'��0�ށ�D/T Q�B��М��D � � �@�й��ҥ@���������Ѐ1�@�@⨐���Y R��Y��A�	@�
@�@�@�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�?D�?�3�4 ��2�4��Y�Y �4
�4�4����4�(O :OLO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�N�`�r������� ��̏ޏ����&�8� J�\�n���������ȟ ڟ����"�4�F�P� $Or���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �f������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o��o�o�a�$PGT�RACELEN � �a  ����`��f_�UP ���e�q'pq p��a_CFG �Fu	s�a0q�Lt��ceqxc}  ��qu4rDEFS_PD �?|�a�p��`H_CONFIG �u�s �`�`d��t��b �a�qP��tcq��`��`I�N7pTRL �d?}_q8�u�PE�u;��w�qLt��qqv�`LID8s��?}	v�LLB 1}��y ���B�pB4Ńqv ��އ؏	�s �<< �a?� �'���A�o�U�w� ������۟��ӟ��#�	�+�Y�v�񂍯�� ��ï
��������/�~u�GRP 1ƪ���a@�j���hs�aA�
�D�� D@� �Cŀ @�٭�^�t������q�p����.� ���Ⱦ´���ʻB�)�	����?�)�c��a>��>�,��Ϻ������ =49X=H�9��
����@�+� d�O���s߬�o߼�����  Dz���`
��8���H�n�Y�� }�������������@4��X�C�|���)���
V7.10b�eta1Xv �A������!������?!G�>¿�\=y�#��{�33A!��@���͵��8wA���@� A�"s�@Ls���� ��"�4FXLsApLr�y�ā��_��@l��@�33q��`s��k��A�nff�a������)�x�� �ar�T�n�t�����	t�KNO?W_M  |uGv�z�SV ��z�r�&����>�/�/G/�a��y�M�M���{ ���	�^r�` (l�+/�/',�$@�XLs����@ ���%�"4�.N�z�+MRM��|-TU��y�c?u;eOADB�ANFWD~x�S�TM�1 1�y��4Garrwa_B�2Sema��?~s�;Co�2���O�7�3An�tena_Full @��VODe� qH��^OpO�O�O�O�O �O�O!_ __W_6_H_@�_l_~_�_�b�72�<��!4�_  �<�_�_N�3�_�_
oo��749oKo]ooo�75 �o�o�o�o�76�o�o�772DVh��78�����7M�A�0��swwO�VLD  �{��/a�2PARNUM  �;]��u��SCH*� 8�
�����ω�3�UPD���[�ܵ+�wu_CM�P_r -��0�'��5C�ER_CHKQ����1�"e�N��`�RS>0�?G�_M�O�?_��#u_R�ES_G�0��{
 Ϳ@�3�d�W���{� �������կ���*� ����P��O� �8`l�������`�� ʿϿ��`�	��� 1p)�H�M���phχπ����p�������V� 1��5�1�!@�`y�ŒTHR_�INR>0/�Z"�5d�:�MASSG� Z�[�MNF�y�MON�_QUEUE a��5�6Ӑ~  #tNH�U��N�ֲ����END�����EX1E�����BE����>��OPTIO�������PROGRAM7 %��%��������TASK_I�,�>�OCFG �ά�]�����DAT�Au#��������2 �O
=�TE�U��^�p������:�  �����=����������4 �� ~� ~ � /xAS�INFOu#� ���Ԕ$��� ���
.@R dv��������/as x� � �;���ȀK_��q���S&ENB-�Hb-&q�&2�/�(G���2�b+ X,{		��=����/O��@��P4$�0���99)�N'_EDIT ���W?i?>��WERFL�-���3RGADJ ��F:A�  �5?@Ӑ�5Wј6��]!֐���?� ' Bz�WӐ<1Ӑn&%�%O�8;��50!�2��7�	H��l�0�,�BP�0��@�0�M*z�@/�B **:�B��O�F�O2��D��A �ЎO�@O	_,X��%�:��H�q��O$_@r_0_�_���Q@WA�� >]�_�_�_o�_o�_ �_
o�o.o�ojodovo �o�o�o�o�o�o\ XB<N�r�� ��4��0���&� ��J������������ �����x�"�t�^� X�j�䟎���ʟğ֟ P���L�6�0�B���f� ��������(�ү$�� ����>���z�t���  Ϫ������l�� h�R�L�^�DX	������0�� ���t$  :�L��o�
ߓߥ��7PREF ��:�0�0
�5IOR�ITYX�M6��1MPDSPV�:n" ��UT��C�6ODU[CT��F:��vNFOG[@_TG�0���J:?�HIBIT�_DO�8��TOE�NT 1�F; �(!AF_IN�E*�����!t�cp���!u�d��8�!ic�m'��N?�XY�3�vF<��1)� �A�����0������� ����' ]D �h������*>��3��9n"OxTf�3>�'��F��G/�LC��4��;LFJAB,  ���F!//%/7/�5�F�Z�w/�/�/�/�3&ENHANCE �2
FBAH+d�?�%;�������Ӓ1�1PORT_NUM+���0���1_C_ARTRE�@��>q�SKSTA*��oSLGS�������C�Unothing?�?O�O�۶0TEMP ��N�"O�E�0_�a_seiban |߅OxߕO�O�O�O�O _�O'__K_6_H_�_ l_�_�_�_�_�_�_�_ #ooGo2okoVo�ozo �o�o�o�o�o�o1 U@e�v�� �������Q��<�u�.IVERSI�	�L��� d?isable'2*KSAVE �N��	2670H7K71|�h��!�/0��9�:� 	^�4�$�ϐ����e��͟ߟ�����9�D�tC-Å_y� 1������ő�����Ǻ�URGE� B��r�WFϠ��-��9�W����l:W�RUP_DELA�Y �=n�WR_HOT %���7��/p��R_NORMALO�V�_�����SEMI���������QSKIPo��97��xf�=�b�a�s� ��H��ʹ��ø����� ���&��J�\�n�4� Fߤߒ������߲�� �� �F�X�j�0��|� �����������0� B�T��x�f�������|��ãRBTIF��5���CVTMOUڞ7�5���DC�Ro��� ��T�B׾�C��1bCӏ&?���q>���=�[H������8��^�������*[F�0�K�HϘ�� <
6�b<߈;܍��>u.�>*��<��ǪP0���2DVh z��������,GRDIO_TYPE  v��/�ED� T_CFGg ��-�BH]��EP)�2��+ �C�u �/�*� �/�?�/%?=�/V? �}?�Ϟ?���?�?�? �?�?O
O@O*Gl?qO ��8O�O�O�O�O�O�O �O�O_<_^Oc_�O�_ _�_�_�_�_�_o�_ &oH_Mol_o�oo�o �o�o�o�o�o�o"Do Iho*j��� ����.3�E�� f� ���x�������� ҏ�*�/�N��b�P� ��t�����Ο��ޟ��:�+���R'INT �2�R��!�1G;� i�{��"���8f�0 ��ӫ�� ����M�;�q�W� ������˿���տ� %��I�7�m��eϣ� ���ϵ�������!�� E�3�i�{�aߟߍ��� ����������A����EFPOS1 1��!)  x ���n#��������� �����/��S���w� ���6�����l����� ��=O����6� ��V�z�  9�]���� Rd���#/�G/ �k//h/�/</�/`/ �/�/??�/�/?g? R?�?&?�?J?�?n?�? 	O�?-O�?QO�?uO�O "O4OnO�O�O�O�O_ �O;_�O8_q__�_0_ �_T_�_�_�_�_�_7o "o[o�_oo�o>o�o �oto�o�o!�oEW �o>���^� ����A��e� � ��$�����Z�l���� �+�ƏO��s��p� ��D�͟h�񟌟�'� ԟ�o�Z���.��� R�ۯv�د���5�Я Y���}���*�<�v�׿ ¿����Ϻ�C�޿@�xy��e�2 1�q� �-�g�����	��-� ��Q���N߇�"߫�F� ��j��ߎߠ߲���M� 8�q���0��T�� ������7���[��� ��T�������t��� ��!��W��{ �:�^p�� A�e �$� �Z�~/�+/� ��$/�/p/�/D/�/ h/�/�/�/'?�/K?�/ o?
?�?.?@?R?�?�? �?O�?5O�?YO�?VO �O*O�ONO�OrO�O�O �O�O�OU_@_y__�_ 8_�_\_�_�_�_o�_ ?o�_co�_o"o\o�o �o�o|o�o)�o& _�o��B�f x��%��I��m� ���,���Ǐb�돆� ���3�Ώ���,��� x���L�՟p������� /�ʟS��w��������3 1��H�Z� �����6�<�Z���~� �{���O�ؿs�����  ϻ�Ϳ߿�z�eϞ� 9���]��ρ���߷� @���d��ψ�#�5�G� ��������*���N� ��K����C���g� �������J�5�n� 	���-���Q������� ��4��X�� Q���q�� �T�x�7 �[m�//>/ �b/��/!/�/�/W/ �/{/?�/(?�/�/�/ !?�?m?�?A?�?e?�? �?�?$O�?HO�?lOO �O+O=OOO�O�O�O_ �O2_�OV_�OS_�_'_ �_K_�_o_�_�_�_�_ �_Ro=ovoo�o5o�o Yo�o�o�o�o<�o `�oY��� y��&��#�\��������?�ȏ����4 1�˯u�����?� *�c�i���"���F��� �|����)�ğM�� ���F�����˯f�� ������I��m�� ��,���P�b�t���� ��3�οW��{��x� ��L���p��ϔ�߸� �����w�bߛ�6߿� Z���~�����=��� a��߅� �2�D�~��� �����'���K���H� �����@���d����� ������G2k� *�N���� 1�U�N� ��n��/�/ Q/�u//�/4/�/X/ j/|/�/??;?�/_? �/�??�?�?T?�?x? O�?%O�?�?�?OO jO�O>O�ObO�O�O�O !_�OE_�Oi__�_(_ :_L_�_�_�_o�_/o �_So�_Po�o$o�oHo��olo�oۏ�5 1����o�o�olW� �o�O�s��� 2��V��z��'�9� s�ԏ���������@� ۏ=�v����5���Y� �}�����۟<�'�`� �������C���ޯy� ���&���J����	� C�����ȿc�쿇�� ���F��j�ώ�)� ��M�_�qϫ����0� ��T���x��u߮�I� ��m��ߑ������� �t�_��3��W��� {������:���^��� ���/�A�{�����  ��$��H��E~ �=�a���� �D/h�'� K���
/�./� R/��/K/�/�/�/ k/�/�/?�/?N?�/ r??�?1?�?U?g?y? �?O�?8O�?\O�?�O O}O�OQO�OuO�O�Ox"_t6 1�% �O�O_�_�_�_�O�_ |_o�_o;o�__o�_ �oo�oBoTofo�o �o%�oI�omj �>�b���� ���i�T���(��� L�Տp�ҏ���/�ʏ S��w��$�6�p�џ ���������=�؟:� s����2���V�߯z� ����د9�$�]����� ���@���ۿv����� #Ͼ�G�����@ϡ� ����`��τ�ߨ�
� C���g�ߋ�&߯�J� \�nߨ�	���-���Q� ��u��r��F���j� �����������q� \���0���T���x��� ��7��[�� ,>x����! �E�B{�: �^�����A/ ,/e/ /�/$/�/H/�/ �/~/?�/+?�/O?5_GT7 1�R_�/? H?�?�?�?�/O�?2O �?/OhOO�O'O�OKO �OoO�O�O�O.__R_ �Ov__�_5_�_�_k_ �_�_o�_<o�_�_�_ 5o�o�o�oUo�oyo �o�o8�o\�o� �?Qc���"� �F��j��g���;� ď_�菃������ˏ �f�Q���%���I�ҟ m�ϟ���,�ǟP�� t��!�3�m�ί��� �����:�կ7�p�� ��/���S�ܿw����� տ6�!�Z���~�Ϣ� =ϟ���s��ϗ� ߻� D������=ߞ߉��� ]��߁�
���@��� d��߈�#��G�Y�k� �����*���N���r� �o���C���g����� ������nY� -�Q�u���4�X�|b?t48 1�?);u� �/;/�_/�\/ �/0/�/T/�/x/?�/ �/�/�/[?F???�? >?�?b?�?�?�?!O�? EO�?iOOO(ObO�O �O�O�O_�O/_�O,_ e_ _�_$_�_H_�_l_ ~_�_�_+ooOo�_so o�o2o�o�oho�o�o �o9�o�o�o2� ~�R�v��� 5��Y��}����<� N�`���������C� ޏg��d���8���\� 埀�	�����ȟ�c� N���"���F�ϯj�̯ ���)�įM��q�� �0�j�˿��ￊ�� ��7�ҿ4�m�ϑ�,� ��P���tφϘ���3� �W���{�ߟ�:ߜ� ��p��ߔ���A��� �� �:����Z��� ~�����=���a������ �����MAS�K 1����������XNO  ����� MOTE�    N_?CFG �Y�����PL_RAN�GUP���OW_ER ��� ��A��*SYS�TEM*P�V9.�3044 �1/�9/2020 �A �g ���R�ESTART_T�   , $�FLAG� $D�SB_SIGNA�L� $UP_�CND4��RS�232r �� $COMME�NT $D�EVICEUSE�4PEEC$PA�RITY4OPB�ITS4FLOW�CONTRO3T�IMEOUe6C�U�M4AUXT���5INTERF{ACsTATU��KCH� t $OL�D_yC_SW �'FREEFR�OMSIZ �A�RGET_DIR� 	$UPD�T_MAP"� T�SK_ENB"E�XP:*#!jFA�UL EV!�R�V_DATA�_  $n E��   	$VAL�U�! 	j&GR�P_   �{!A  2 ��SCR	�� �$ITP_��" $NUMΞ OUP� �#TO�T_AX��#DS}P�&JOGLI�FINE_PCdn�OND�%$�UM�K5 _MIiR1!4PP TN?8�APL"G0_EX�b0<$�!� 814�!P=Gw6BRKH�;&{NC� IS �  �2TYP� �2�"�P+ Ds�#;0BS�OC�&R N�5DU�MMY164�"S�V_CODE_O�P�SFSPD_�OVRD�2^L�DB3ORGTP; LEFF�0<G� �OV5SFTJRUNWC!SFpF5%3oUFRA�JTO��LCHDLY7R�ECOVD'� WaS* �0�E0RO���10_p@  � @��S NVE�RT"OFS�@C� "FWD8A�D4A��1ENABZ6�0T�R3$1_`1FD}O[6MB_CM�!zFPB� BL_M��(!2hRnQ2xCV�"�' } �#PBGiW|8A�Mz3\P��U�B�__�M�P�M� �1�AT�$CA� �PD�2��PHBK+!:&aI�O�4 eIDX+bPPAj?a$iOd�7e�U7a�CDVC_DBG"�a;!&�`��B5�e1�j�S�e3��f�@ATIO� ���AU�c� �S�AB
0Y.#0�D���X!� _�:&S�UBCPU%0S�IN_RS�T, 1�N|�S�T!�1$HW_C1�"]q.`�v��Q$AT! � �_$UNIT�4�p>�pATTRI= �r�0CYCL3NE�CA�bL3FLTR_2_FI9a7�c�,!LP;CHK�_�SCT>3F_ƥwF_�|8��zFS8+�R�rCHAGp�py��R�x�RSD�@`'�1E#&7`_T�X�PRO�`@S�EMOPER_0�3Tf��]p� f��P�DI�AG;%RAILAiC�c4rM� LO�04�A�65�"PS�"�2� -`�e�SPR�`S&.  �W�Ctaf�	�CFUNC�2~�RINS_T.!`(�w��� S_� ��0�P�� 	d��W�ARL0bCBLCUR��єAʛ�q͘ƘDA�0���ѓʕLD @,a3��!��8�3�TID�S��!�� $CE_RIYA !5AFDpPC�~��@��T2 �C�9#�b{QOI�pCVDF_LE��#0(!��LM�SFA�@HRgDYOL1	PRG8��H��>1(�ҥMUGLSE =#Sw3��$JJJ6BKGFK�FAN_ALML�V3R�WRNY�HGARD�0+&_P "B��2Q���!�5_�@�:&AU�Rk��TO_SBRvb��� �ƺ�pvc�޳MPINF�@�q�)���'REG'd~0V) 0R<�C�1DAL_ \2sFL�u�2$MԐ (�#S��P� `�gśCMt`NF�qsO!NIP�q5P��IPP� 9a$Y��! �"�!�� �o3EG0P��#@��AR� �c��52�����|5AX�E�'ROB�*REMD�&WR�@�1_=݆�3SY�0ѥ0_�S�i�WRI�@�ƅpST�#��0*@� �q!	���3��� B� �At��3�D�POTO�9� �@ARY�#��0!��d�!1FI�0��$LINK��GkTH�B T_����A��6�"/�XY�Z+"9�7G�OFF��@�.�"���B� l����A3$ ��FI�p���4�4l��$_Jd�"(B�,a������8�"q�������Ck6DUtR��94�TURT�!XZ�N����Xx��P��FL/�@s��l��P��30�"Q +1� K
0M:$�5�3]q7�SuD�Sw#ORQɆ�!�����Q7�
�0O[�ND�=#�!�#�1OVE8��M ���R��R��Q�!P.!P! OAN }q	�R����990�  �brJ9V����Lv�!ER1��	8�!E�@n D�A��p�嘕Ă���v�AX�C�"��`�q� s���0~3� ~F�~e�~�~E�~1��~Ҡ{Ҡ� Ҡ�Ҡ�Ҡ�Ҡ� Ҡ�Ҡ�Ҡ�!)oDEBU}s$x�`��삼!R*�AB��a8A2V`|r 
�"�c���%�Q7� 7�173�7F�7e� 7�7E�����.��LAB����yp��cGRO�p��}��PB_ҁ ��1C���ð�6�1���5���6AND��8p�a3���-G �Q����AH�PH�p2�NTd��Cs@VEL؁�}A��F?�SERVEs@��� $����A!�!�@POR}�KP��b�A�B���	���$�BTRQ�
��CH��@
�G��2	��Eb��_  qlb��Q�ERR��RI�P�@�FQTO	Q�� L�}��YV�ĀG�E%�\���CRE�  �,�A�EP
�RA~�Q 2 d�R�7c��T�@ ��$F ׂ��m����BOC��P � 8[COUNT��ќ��SFZN_wCFG�A 4�p%��rT\zs�a�#`p�Jp c%d�� �� MGp+����`�OGp�eFAq����cX8еk�ioQ��'ѴD�p8�Pz���HE�LA�-b }5��B_BAS\�RSR$�`�2�SH��L�!p1�W!p2DzU3Dz4Dz5Dz6Dz�7Dz8�WqROO0���P�1�NL�� ��AB�C
�"pACK��&IN�PT+�W�Up��	�k��y_PU8�,~�|�OU�CP��%��s�Vl���YTPF?WD_KARKQ-�&:PRE�D�P����QUE$�Ā9 )���~���IU��#s/�p��@�/�SEM1�ǆ1�A�aSTYf�tSO����DI�q���Qc��X��_TM>9�MANRQ �/��END��$KEYSWITCH2��G����HE)�BE�ATMz�PE��L�EJR���0x�UF�F���G�S�DO_H�OM��Oz��pEFPR��SbJі��u�C��O��7P�QOV�_M��}�c�IOC�M���1�BsHK�� D,�&�a`	U2R��M��a�r +��FORC*�WARn���� uOM��  @�$�㰰U��P�1��g���e3��4�1.��S�P�OW�Lz��R%�U�NLO�0T�E�D��  �SNuP��S.b 0N��ADDa`z�$S{IZ*�$VA�0~�UMULTIP�r�P���Az� � $��ƒ����SQc�1CFPv�F'RIFr�PSw����ʔf�NF#�ODBUx�R@w������F��:�IAh�����������S"p�� �  �cRTE���SGL.�T�x�&�C`Gõ3a�/�STM�T��`�P����BW<9 0�SHOWh�q7BANt�TPo���@E�����PV�_Gsb �$PaC�0�PoFBv�-P��SP��A�p����PVD��rbw� �+QA002D .ҝ�6ק�6ױ�6׻��6�54�64�74�8*4�94�A4�B4و� 6ׇ17�}�6�F4�  ��@�����Z����t�U1��1��1��1��U1��1��1��1��U1��1��23�2@�U2M�2Z�2g�2t�U2��2��2��2��U2��2��2��2��2��2��33�����M�3Z�3g�3t�3���3��3��3��3���3��3��3��3���3��43�4@�4�M�4Z�4g�4t�4���4��4��4��4���4��4��4��4���4��53�5@�5�M�5Z�5g�5t�5���5��5��5��5���5��5��5��5���5��63�6@�6�M�6Z�6g�6t�6���6��6��6��6���6��6��6��6���6��73�7@�7�M�7Z�7g�7t�7���7��7��7��7���7��7��7��7���7��hbVPv�U�B �@�09r�
o�V���A x� �0R���  ��BM�@RP�`�4Q_�PR�@[U�AR��D�SMC��E2F_�U��=A ��YSL|�P�@ �  � ֲ>g�������iD��VALU>e�pL��A�HFZAID_L����EHI�JIh�$FILE_ ��D�dc$Ǔ�PXCSA�Q� h�0!PE_BLCKz�.RI�7XD_CPUGY!�GY��Ic�O
TUB���R�  � PaW`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q��TJ��U�Q�T�Q�UH`��T`�T@�T2L��_LIz�  ]�pG_OT�P_EDIU�-b�`7c ?bة�pBQh�~�� �TBC2 �! �%�>��P���a�7aFTτ�d݃T�DC�PA�N`�`M0�0�f�a�gTH��U��d�3�gR�q�9�ERVEЃt݃t�	��a�p�` "�X -$EqLE�NЃRt݃Ep�pRA�v��Y@W_AtS14Eq�D2�wMO?Q�	S���pI�.B�A�y��4Ep�{DE�u��LgACE �CCC�.B��_MA��v��w�TCV�:��wT,�;�Z�P���sѨ~��s�J�A�MD����J���uā
�uQq2ѐ���݁l�s�JK��VK�� ����	���J�����JJ�JJ�AAL�<��<�6��2:�5�cm�N1a�m�(,��DL�p_\�Q�0ApCF
�# `�0GROU�@J�Բ���N�`C^�ȐRE�QUIRrÀEBqUu�Aq��$T�p2"��Bp薋a	��d�$ \?@qhAPPmR��CLB
$H`�N;�CLO}`K�S��e`��u
�aI�% �3�M�`�l��'_MG񱥠C �"Pp����&���BRK���NOLD����RTCMO6a�ޭ��J6`�P>��p��p��pPZ��pc��p6+�7+��<����e&� �lr��������PATH���������qx�����%0A��S�CAub��<���INFDrUC�p�q�C�KUM�Y�psP�� ��A q/ʤ�/�E�/��PAYLOA�J{2L�0R_AN�ap�L�Pz�v�jɆ����R_F2LSHRt��LO{�R����|���ACRL_�q �����b�d�H�@B�$H��"�FLE�X>�$�`J�f' P(��o�o+�p�>�Du( : Qcv�p����fe��po��|F1���-瀢�����]�E ��*�<�N�`�r��� ��4�Q�������A�c� ��ɏۏ���T��2�X:A������ ����)�;�?�H�6��Z�c�u�����.`BJ��) ��`��˟ݟ��`�0ATF�𑢀E�L��(a��J�(v��JE۠CTR���A�TN�1�HA_ND_VBB>�ܯ@�* $��F24���d�CSW>�=s���+� $$M �����0ˡ�ڡ������A�@g����AD)��A���@˪A٫AA� ��`P˪D٫�D�PȰG�P�)S�Tͧ�!ک�!N�DY�P9����#%��Fp ���Ѫ���i����������P3�<�E�N�W��`�i�r���J�e,1 ��ԓ� n�5<m��1ASYMص.@	�ض+A������_`��	���D� &�8�J�\�n�Ju�&���ʧC�I��S�_VI�o�Hm��@V_UANVb�@
S+��J� "RP5"R��&T��3TWV �͢���&��ߪU��a/�7�w��`HR`�ta-��QQ�1�D)I��O�T����PN��. ; *"IAA*���$aG�2C2cJ��$��I��P / �� �ME��� Mb�R4AT�PPT@�@� ��ua���PАl@zh�a�iT�@��� $DUMMY}1E�$PS_D�RF�w�$�fn3�FLA��YP����b}c$GLB_T��Uuu`1�� ��EQa0 X(����ST����SBR��PM21_V��T�$SV_ER��O�_@KscsCLpKrA���O'b�PGL�@E�W��1 4��a+$Y|Z|W�s����AN`�  ��sU�u2 ��N��p�@$GIU{}$�q 1�t�p��3 L���v^B�}$F^BE�vNE+AR��NK�F8����TANCK�  ��JOG��� �4� $JOIN�T�����uMSET.��5  �wE�H�� S����� ��6��  MU��?����LOCK_F�O����PBGLV�HGL�TEST�_XM>���EMP�t����r̀$1U�Гr��22���sB,�3���Ҁ,�1Mq�CE���sM� $K�AR��M�STPD�RA�pj�a�VECX��{�e�IU,�41�{HEԀTOOL�ڠ�V�RE��IS�3����6N�A�AC)H���5��O�}cj�d3���pSI.��  @$RAI�L_BOXE���ppROBO��?�~pqHOWWAR*�x��`�ROLM�b B���S��
�5����O_F� !ppHOTML5�Q�����AP�QGU�C�H��7m�
��R
��O��8m��v�z��!p�sOU��9 	tpp(�14A�̀���PO֡%PIP��N��
�ڑS��,�����CORDEaDҀް̠5�XT���q)���P� O4` �: D pOBP!"Ҁ{�j��cp�j�^@$SYSj�A�DR#�Pu`TCH�� ; ,��E�N�RZ�Aف_�t�״�>��PVWV�APa< � �p��r�UPREV_�RT]1$EDI}T�VSHWR��7v;���q�@D�_`#R�+$H�EADoA�Pl�A�$�KE�q�`CPS�PD��JMP��Ld�U� R��d=r�TO�϶I�S#Ci�NE��$_TIC�K�AMX�AS���HN-q> @pt������_GP֜�[�STYѲ�LAOq���Ҩ�?�5
�Gݵ%$���tu=7pS !$Q ��da�e!`�fP�0ևSQUd� ��b�ATGERCy`|�pS�@ �pCp����d�%Oz`mcO�IZ�d�q�e�aP�RM��a8����PU�QH�_DO=�ְXuS��K�VAXIg�f�1�UR� ��$ #�Е��� _�����ET��Pۂ���5�f�F�7g�A�!�1U�d9�2;]��TSR|Al �о���#��5�� #��#�)#�)i�>' i�N'i�^&{����){�H���2��C����C���WOiO{O�D�qSSC�p B hppD1S(�a�`SP`�ATL �I����~�bADDRES��=B'�SHIF��"��_2CH#��I\&p��TU&pI�� C͢CUST}O��AC�TV��IbDȲ,��0�
�
��U�R`E \�����f�7���tC�#	���F���irt�TXSCR�EEl�F�P��T�INA�s�p��tpb����0G T�� fp,⧱eqBp&uᦲ8u�$#�RRO'0R�`��}�!Ce�pUE��GH ��0���`S�qN��RSM�k�UV�0���V~!�PS_�s�&@C�!�)�'C��Cǂ�z"� 2G�0U�E�4Ibvr�&8�G+MTjPLDQ��Rp��z�BBL_�W��`R`J �f�>2O�qJ2LE�U3"��T4RIGH^3B�RDxt�CKGRĦ`�5TW��7�1WIDTH�H����a�a����UIu�E9Y��QaK d�p���A�J�
�4�BAC�KH��b�5|qX`F�OD�GLABS�?�(X`I�˂$UAR(�9@��0^`H4!� L 8�QR�_k��\B_`R�p͂�����HBO�R`M���w0Uj0�CRۂM�LUM�C��� �ERV�\!I�PN�E�4NV`��GE`=B#���]�t�LP�E��E��Z)Wj'XPz'XԐ&Y5$[6$[7$[8	R���3�<����fԑŁS���M�1USR�tO <��^`U�r�rsFO
�rPRI���m����PTRIP��m�UNDO��P�p��`m�4�l�C�#���� �QWB�P7�G �s�Tf�H�RbOS�agfR��:">c��.qR��s�~�b*��!$�	UQ.qS�o�o�#R�)�>cOFF���pT� �cOp 1�R�t/tS�GU��P.q��JsETw�1�SUB*� f�E/_EXE��V��>c�WO>� U�`�^g��WA'��P�qz!@� V_DB�s��p�2SRT�`
�V0�Q�r��OR��u'RAU��tT�ͷr�q_���W |%��͸OWNA`޴$GSRCE � ��D��<\��MPFIA�p��ESPD����� �C���Gƒ�@+�5��!GX `�`�r޴�n��COP�a$��C`_w������rCT�3�q���qƒp���@� Y"SHADOW�ઓ@�?_UNSCA��@���4M�DGDߑ��E�GAC�,Me�G��Z (0NOX�@�D<�PE�B��VW�S�G���![o � ��VEE#��ڒANG�$��c�薴cڒLIM_X �c��c� ����#`��`� 퐾�VF� ��s�VCCjв�\ՒC{�RAlצ���\RpNFA��Z%�E��Z`G� f^0[�C`DEĒ��� STEQ1���@ �ꁻ@I��`+0���p�`����P_A6��r���K��!]�# 1Ҡ�����\�ȫсCPC�@]�DRIܐ\�͑V#Ѐ����D�TMY_UBY�T���c��F!���bY�븲���P_V��y��LN�BMQ1�$��DEY��EXX�e��MU��X�M� US�!���P_AR����P� ߖG��PACIr�ʐf�ᔀ���c�´c���#�EqB��a.2B���Ч^ ܀GΐP����)�D�R~``�_ �0�@3!�1zr	�e�R�SW��p�00��$S�6�O�Q�1A� XӚ#�E�UE��00���C�HKJ�`�@�p���U� �EA�N�ٖp�pX��MR�CV�!a ��@O*��M�pC�	��s����REF*7
��� �����/��P��@��� @��b��֗�_Y��� ���ۣ��Q$3���8��?��$b �����%���Q��$GROU� �c�����ʠ]��I2^0��U` 0_�I,�o V� ULա`��C&�frAaB�?�NT�� �������A���Q��K�L����õ��A���Qr��T a$c t�`3MD�p8�HU���vSA�CMPE �F  _�R r�p@����XS	���GF/�b#d, �&�@M�P^0۰UF�_C !���z �RO h0"+���@���0C��UREB���RI��
IN�p������d��d��ca�IN"E�H�y��0V�a-�걗�3�W����`���C��i�LO��}�z�@0�!�QNSI��݁���c$&�c$&^.�X_PE-YW+'Z_M�ڒW�Iӑ$�" �+R�'rR;SLre �/�IM
`�RE�C7�Gd�۰�̵ҭ�q��� �u��Ȑ���`���S_P�VnP *��IA�vf �~pHkDR�p�pJO�P���$Z_U�P��a_LOW��5�1J�dA��LINubEP?�tc_i�1�1���@�G1@��V��xg 5X�P�ATHP X�CACH$�]E��yI��A��{�C)�ID3F�A�ETD�H��$H�O�pղb@�{��d6�F�����p�PA3GE�䁀VP�°��(R_SIZ��2TZ�3�-X�0U�q�MP\RZ��IMG���sAD�Y�MRE���R7WGP��8�p��ASYNBUF�VRTD�U�T7Q�LE_2D-��U�J�`CҡU1��Qu���UECCU��VE�M��]EDb�GVIR�C�Q�U�S�B�Q�L�A��p�NFOUN^_�DIAG�YRE�GXYZ�cE�W� �h8�dpqa`T��2IM�a�V|be��EG/RABB��Y�aЗLERj�C4���FC-A�6504x��7u��� BE��h'�>`�CKLAS_@l�8BA��N@i  G��IT��� @ݲմ$BAƠwj �!q�eb��uTYSp�H����2B��I�t:b�f��B)�gEVE����PK��؂fx��GI�pNOt��2�\r_HO��>��k � ���
8�Pi�S�0ޗ���RO�ACCEL�?0=���VR_�U�7@�`��2�p��ARF��PA��̎K�D���REM_But M�rJMX �l�t>�$SSC�Uk� #���QN@m �� �S�P�NS����VLEX�vn =T�ENAB 2¼W@��FLDRߨF�I�P�t�ߨ(Ğ���2P2HFo� ���V
Q MV_PI��8T@�H���F@�Z� +�#��8�8#��sGAB���LOO󣎔�JCBx��w"SC�ON(P�PLANۀ�Dp�3F�d�v�9PէM��Q ;����SM0E�ɥ�8ɥWb 72$`<�8T��,`�RKh"ǁVANC���@AR_Ou N@p (�-#<#c��c�2 w�A/�N@q 4������`	�^�� w�N@r hn���1�^�&OFF`|�p��`��`�DEA�
��P,`SK�DMP6V{IE��2q w���@���rs < {���4���r{7���D��Ȭ!CUS�T�U��t $�G�TIT1$sPR\��OPTap� ��VSF�йsuB�p�0`r&��1SMOwvI�|�ĄYJ�����eQ_WB��wI���� @O3��@�XVRxx�mr��T��
�Z�ABC��y �op����)�
}qZD�$�CSCH��z Lu����`�2�%PC ��7PGN ��<�<�A��_FUNH��@�)P�ZIPw{,I��LV,SL��~�}��ZMPCF���|��E����X�DMY_LNH�=�C�� ~��} $�A�� ]�CMCM� C�,SC&!��P�� �$J���D Q�������������a_�Q,2����UX�a>\�UXEUL��a ������(�:�(�J���FTFL��w�7�Z�~Zp+�T6����Y@Dp�  8 $�R�PU��> EIGH����?(�iֱ�q�0��et� �a�����$B�0�0@�}	�_SHIFD3�-�RVV`Fcв�		$5��C�0��&!������b
�sx�uMD�TR��V̱���SPH���!�� ,������� ��4A�RYP��%������%��"��%!  �H�(UN0���"�2 �����ɐ�q0�GSPDak����P��O�����0��첱��"!NGVER`q �iw+I�_AIRPURG�E  i  �i/�F`E�Tb� ��+1h2ISOLWC  �,�"!�%��P+��_/*OB��Dm�?�@�!H?771  34n?��?�9� `�E/#�)x�� S232�� 1�i� L�TEk@ PEND�A�341 1D�3<*? M�aintenance Cons B��? F"O,DNo UseMJOO�nO�O�O�O�O2�2N�PO;� 19%v�1CH=� �.��		9Q_!�UD1:___RS?MAVAIL/�/%��A!SR  ��+��H�_�P1�T7VAL.&���P�(.�YVL�}� 2|i�� D��P 	�/_oUQNo�o rci�o�g�o�o�o�o �o*,>tb �������� �:�(�^�L���p��� ����܏ʏ ��$�� H�6�X�~�l�����Ɵ ���؟�����D�2� h�V���z�������� ԯ
���.��R�@�b� d�v�����п����⿀��(�N�<�r�i��$SAF_DO_PULS. jQp�����CA� �/%��&0SCR ��`X���0�0
	14�1IAIE���b vo$�6�H�Z� l�~�ߢߴ������߬���HS��2�%�����d1�(�8�8rb��� @�"k� }���T�h� J`���_ @��T7 �����#�0�T D��0�Y�k� }��������������� 1CUgy�O<�Ef������  �5;�#o�� 1p�U��
�t��Di��������
  � ��*������gy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7O<A���`OrO�O�O�O�O �O�O�O?O�_._@_ R_d_v_�_�_�_�_�Q _�R0MJTo !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ JO��'�9�K�]�o� ������_ɟ۟��� �#�5�G�Y��_�U�_ �ҙ�����ϯ��� �)�;�M�_�m����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B�T�f�;�?�q߮� ����������,�>� P�b�t�������������������Y��	123456781�h!B!�)���F����� ������������  ��;M_q�� �����% 7I[l*��� ����//1/C/ U/g/y/�/�/�/n� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? O�/)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_O_�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�op_ �o�o�o/AS ew������ ���o+�=�O�a�s� ��������͏ߏ�� �'�9�K�]������ ����ɟ۟����#� 5�G�Y�k�}�������"��s�կ�w����0�L�CH  �Bpw�   ��=�2�� }� =�
���  	�o�ί���ǿٿ���r���� ��@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖ�%Ϻ��� ������&�8�J�\� n����������� ���"�Q�*������;�<M���D���  �]�w�*��Z򛱛�t  �d�����*�`*��$�SCR_GRP �1*P�3 � �*�� 6�	 �� 
��<�+*�'pUC|@��y�yD� W�!��y�	M-10�iA/7L 12�34567890ڙ�� 8��M1T� � �
�	L���	Č� N 
���Y���y�
M_	P������ ,��#H�
 ���1/�@A/g/y/H�ߙ! T/�/P/�/3��+���/B�S��,?*2C4r&Ad�R?  @s�j5N?�7?��7&2R���?}:&F@ F�`�2�?�/�?�?O O-OSO>OwObO�O=�j1�2�O�O�O�O�DB��O�O;_&___J_�_ n_�_�_�_�_�_o�_ %o�5j�eSgxo6����uo�o�b�1�B̃|3�oh0�4j9j9B� w�$Y̯@HtA�Nhcu�/�%Ipp�drsq ����z�q�x� �.� (&�*�2� D�V�oz�e��������ECLVL  Ψ���iqpQ@���L_DEFAU�LT ���s�փHOT�STR�qq��MIPOWERF���H���WFDO�� �RVENT 1ɁɁ�� L!DUM�_EIP�����j�!AF_INEx‧���!FT}��֞����!-/� ���F�!RP?C_MAING�)�q�5���Y�VISb��t����ޯ!TP&ѠPUկ��dͯ*��!
PMON_POROXY+���e��v��D���fe�¿!�RDM_SRV�ÿ��g���!R�,*ϑ�h��Z�!
�[�M����iIϦ�!RLSYNC�����8����!R3OS|���4��>��!
CE�MTC�OM?ߓ�k-ߊ�!=	S�CONS�ߒ��ly���!S�WA'SRCݿ��m��"�;!S�USB#�n�n�!STMC��o]����� ѳ����,���P�V��ICE_KL ?�%d� (%S?VCPRG1S�����2�������o����4������5��6;@��7ch��H���9���� %��������0 ����X�����- ���U���}��� � /���H/���p/ ���/��F�/��n �/��?��8?�� �`?��/�?��6/�? ��^/�?��/X�j�� q���#OhO��lO�O{O �O�O�O�O�O�O _2_ _V_A_z_e_�_�_�_ �_�_�_�_oo@o+o doOo�o�o�o�o�o�o �o�o*<`K �o������ �&��J�5�n�Y����}���ȏ���^�_D�EV d���MC:�4����GRP 2�d�
@�bx 	�� 
 ,V�
@�s�Z������� �����ߟ��@� '�9�v�]�������ЯP����۫Y�
@
@�ܯ
@1�4�]� ��j�����˿Ӵ��� ����0��T�;�M� ��qϮ��[�!��ϡ� �ߡ�K�!�^�p�� ��s�Y��ߩ�����
���@�'�d�v�� y��^���������� %��I�0�Y��f��� �������������3��T7]�e��� �z�����1 Ag"�r�� �=������ !/G/���R/�/�/�/ �/�/"�/�/??C? *?<?y?`?�/�f?�? �?�?�?�?-OOQO8O aO�OnO�O�O�O�O�O _�O)_;_"___�?�_ �_L_�_�_�_�_�_o �_7oo0omoTo�oxo �o�o�o�o�o!x_ E�oU{b��� �����/��S� :�w�^�p�����я��d �X�ZI6� r 	 @�Z��0�+A�����dBjBA�=��������B����AZ.�AĊ��+�A.��Q�B����5�\��i6�A��u��'����%�Ꮛ�%P�EGA_BARR�A_ESTEIR�A����X�T����?=��=X���7
�?�>��A���瓟�����&���������A�xP��f��U�'A�j���´�B�:��<�3�����jB]+�0�T��%�T����d�ʐ���>�pc�?��7�ԳT�@6��A�_���0n�����·�Ak���۸I�K9F�A�G�����B!v,�-���C3�����pBM�>�#�b�(��Y�������HX��?L!���Q��B���AJ���Xk�@fD�3��O�A��������Y�w���.B��B�;��C�H�z�B�?����6���-Ϙ������n��=]����V@���?,����Ö� վ��e�Ak��������OY�A�������AB�J��;%�C$4��aƿBXZ9@���
���ߘ�Ţ��� �ԭ(��^�_��-\¯ԡ�Q�گ���+�������������ߔ�ᶢ���*נ�6��>�ԯb���zװ}
��BM��`s��x�U<�߿�7@6|=�����$�6��� N�@���b�G���L�}�������x7���~K@����V�+A>r��rF��������Y@+�@�<�B��|�A�F�����B)���,o�?ɇ���~0��0~@6�Z� Q�杚��������A�ߍ�]ܖA����������2[����>�ȥA��=��³�NB ��$�w?�dj���to�7\��
�.�%��Z�����A������*�@Ve��B� ������YN�#��BD�	����9A����gB#
q��3��C4#��,?[BVM����COLOCA_PRENS����X�\{B*3Vhz����p���/
&�M�/ (/:/L/^/p&�z/�/�/�/�/�/X�N&�v��*�@�n4�B-N��v�B��������9���z��@�k'@л���آjA������QB!dD���R?�o�^��CU�Z? ?O~?�?uO{B�� �O�O�O�O�O�O�O _ G__x_f_�_�_ �_�_�_&_L_o\_�_ Po>otobo�o�o�o�_ �o"o�o�o&L: p^��o��o�� �� �"�H�6�l�� ���\�Ə���؏� ���D���k���4��� �����ԟ
�L�1� C������d������� ���$�	�H�ү<�*� L�N�`����������  �����8�&�H�J� \ϒ�Կ���������� ���4�"�Dߚ��ϑ� ��j��߲�������� 0�r�W�� ���� ��������J�/�n� ��b�P���t������� ��"�F���:(^ L�p����� � 6$ZH~ ���n�j�/ �2/ /V/�}/�F/ �/�/�/�/�/
?�/.? p/U?�/?�?v?�?�? �?�?�?OH?-Ol?�? `ONO�OrO�O�O�OO 4O_DO�O8_&_\_J_ �_n_�_�O�_
_�_�_ �_o4o"oXoFo|o�_ �o�_lo�o�o�o�o
 0T�o{�oD� ������,�n S�����t�����Ώ ���4��+���ޏ L���p�����ʟ�� 0���$��4�6�H�~� l����ɯ������  ��0�2�D�z����� �j�Կ¿����
� ,ς���yϸ�RϬϚ� �Ͼ������Z�?�~� �r�߂ߨߖ��ߺ� ��2��V���J�8�n� \�~�����
���.� ��"��F�4�j�X�z� ������������� B0f����V xR���> �e�.���� ���/X=/|/ p/^/�/�/�/�/�/�/ 0/?T/�/H?6?l?Z? �?~?�?�/?�?,?�?  OODO2OhOVO�O�? �O�?|O�OxO�O_
_ @_._d_�O�_�OT_�_ �_�_�_�_oo<o~_ co�_,o�o�o�o�o�o �o�oVo;zon \������ ����4�j�X��� |����ُ������ ��0�f�T���̏�� ��z��ҟ����� ,�b�����ȟR����� �ί���j���a� ��:���������ܿʿ  �B�'�f��Z��j� ��~ϴϢ������>� ��2� �V�D�fߌ�z� ������ߠ�
���.� �R�@�b���߯��� x��������*��N� ��u���>�`�:����� ����&h�M�� �n������ @%d�XF|j �����<� 0//T/B/x/f/�/� /�//�/?�/,?? P?>?t?�/�?�/d?�? `?�?O�?(OOLO�? sO�?<O�O�O�O�O�O  _�O$_fOK_�O_~_ l_�_�_�_�_�_�_>_ #ob_�_VoDozoho�o �o�oo�o�o�o�o�o R@vd��o�  ������N� <�r�����b�̏�� ��ޏ ���J���q� ��:�����ȟ���ڟ ��R�x�I���"�|�j� ����į���*��N� دB�ԯR�x�f����� ����&�����>� ,�N�t�bϘ�ڿ���� ��������:�(�J� p߲ϗ���`��߸��� ��� �6�x�]�o�&� H�"���������� P�5�t���h�V�x�z� ��������(�L��� @.dRtv��  �$�<* `Np����� ��//8/&/\/� �/�L/�/H/�/�/�/ ?�/4?v/[?�/$?�? |?�?�?�?�?�?ON? 3Or?�?fOTO�OxO�O �O�O�O&O_JO�O>_ ,_b_P_�_t_�_�O�_ �_�_�_�_o:o(o^o Lo�o�_�o�_ro�o�o �o�o 6$Z�o� �oJ������ �2�tY��"���z� ����ԏ�:�`�1� p�
�d�R���v����� П���6���*���:� `�N���r����ϯ� ����&��6�\�J����¯�����$�SERV_MAI�L  �����ʴOUTPUT�ո�@�ʴRV 2j� � � (r�������=�ʴSAV�E���TOP10� 2� d 6 rƱ���� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t������n�YPY��F�ZN_CFG f��=���J���GRP 2���g� ,B  � A �D;� �B �  B4~=�RB21I�oHELL��f�e�)�*�=�����%RSR��� ���&J5 G�k�������.�  ��/>/P/"\/1��X/1�2��U'&"2��dh,g-�"EHKw 1S �/ �/�/�/#?L?G?Y?k? �?�?�?�?�?�?�?�?�$OO1OCO?OMM� S�ODFT?OV_ENBմ��e��"OW_REG�_UI�O�IMI_OFWDL~@�N��BWAIT�B �)��V��F�YwTIM�E��G_�VA԰_�A_UNcIT�C~Ve�LC�@WTRY�Ge�ʰ�MON_ALIA�S ?e�I%�he��oo&o8oFj�_ io{o�o�oJo�o�o�o �o�o/ASew "������� �+�=��N�s����� ��T�͏ߏ����� 9�K�]�o���,����� ɟ۟ퟘ��#�5�G� �k�}�������^�ׯ �����ʯC�U�g� y���6�����ӿ忐� ���-�?�Q���uχ� �ϫϽ�h������� )���M�_�q߃ߕ�@� �������ߚ��%�7� I�[�������� r������!�3���W� i�{���8��������� ����/ASe �����|� +=�as�� B����/�'/ 9/K/]/o//�/�/�/ �/�/�/�/?#?5?�/ F?k?}?�?�?L?�?�? �?�?O�?1OCOUOgO yO$O�O�O�O�O�O�O 	__-_?_�Oc_u_�_ �_�_V_�_�_�_oo�c�$SMON_�DEFPROG �&���Aa� &*S?YSTEM*obg� $JO0dR�ECALL ?}�Ai ( �}<�copy md:�place_ba�rra_pren�sa.tp vi�rt:\temp�\=>10.10�9.3.62:1?2944 4bo�o��o	w}7�fickup�o�o�c�ofx�~=�esumir?_furad�o<��d���x�f�ss�em_receptor��Z�l�~��#vco-�?�Q������ }:�edr�op*�defeito���oُj�|�z8�.�_15�G�W�0�������_2��ş`ןh�z���_33��E�W����|xy�zrate 61¯4 ��ͯ^�p���:t
�11 C�:� L�ݿ���&���ʿ [�m�ϒ���6�Hω� �����"ϴ�����i��{�{��c8460 :�L������u�tpdisc 0�� ����[�m���wtpconn 0��3�E�W������|6�bfrs:o�rderfil.�dat��mpback�����e�w�
�}-�db:*.*2����K����� v1xF�:\��' �� ��P`r�r2a% 7��Q���̨ ��]o���&s�c?esteir������w;��`���n4���	/k/}/y4 �k2/D/��R/�/�/? ��s,/�/���/j?|? /�o�D?�/�?�?� �?>�?fOxO�� �;O��O�O_'%� �O�OZ_l_~_�O��4_ F_�_�_�_z9�/� �_���_hozo���� EoUo�o�o�o�o/��o �odv���?Q ����߫ܺ�]� o�����5�G���� ���!���ŏ׏h�z� O�1��_U�������������ӟd�v�����$SNPX_AS�G 2������� �XC%���Я  ?����PARAM ����� ��	��PӤ��Ө$������O�FT_KB_CF�G  ӣ����O�PIN_SIM + ���}����������RVNOR�DY_DO  �)�U���QSTP/_DSBi��Ͼ��SR ��� � &#�D�O��O�:�TOP_ON�_ERRʿ��o�P_TN ������A��RIN�G_PRMy�ܲV�CNT_GP 2���!���x 	 ���ϗ��#��Gߔ��VD��RP 1��"�8Ѩ�*߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�}�z����������� ����
C@Rd v������	 *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? [?X?j?|?�?�?�?�? �?�?�?!OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLosopo�o�o �o�o�o�o�o 9 6HZl~��� ����� �2�D��V�`�PRG_CO7UNTJ���{�'ENB��}�M��L����_UPD 1>'�T  
k��� ���"�K�F�X�j��� ������۟֟���#� �0�B�k�f�x����� ����ү������C� >�P�b���������ӿ ο����(�:�c� ^�pςϫϦϸ����� �� ��;�6�H�Z߃� ~ߐߢ���������� � �2�[�V�h�z�� �����������
�3� .�@�R�{�v������� ������*S�N`r���t�_INFO 1��Ҁ� 	 ���3@��1�?�|�?���9 B���ƓA�&����ߌ��I��@L>  A��e ?�" >�a� A�  &Cj��D����3���u�B� ����YSDEBU)G����� dՉ�SP_PASS���B?+LOG ���� � s ��  �с��UD1:\x;$�<"_MPCA-�셽/�/�x!�/ �쁝&SAV �D)��%d!|"�%��(SV�+TEM_TIME 1D'��� 0  -g�#/�()��#�-M7MEMBK  �сd d/�?��?�<X|Ҁ�3 @�?C�O:O�JLOmOzI�J
! %@p1�O�O�O�O "3 __$_6_H_Z_l_ �n_�_�_�_�_�_ �_�_o"o\�e1oVo hozo�o�o�o�o�o�o �o
.@Rdv0���O5SK�0�8����?���F�Ҁ�H2OJ�AJ� ��C�A\O4����(�O"�Oя�b�ݏw_�O �` 9� ��0�9�g�y���
�L����ӟ���	��� $�C�7o g�y���������ӯ� ��	��-�?�Q�c�u�����������T1SVGUNSPD%%� '%��2M�ODE_LIM #a9"ܴ2�	�� D-۵ASK_?OPTION �9�!F�_DI ENB  U�%f��BC2_GRP 2!�u#o2��N���C���ԼBCCF�G #��*< #6�*�`ߐI� 4�Y��jߣߎ��߲� ��������E�0�i� T��x��������� ���/��S�>�w�����t���u�����c� ��	B-f�.� �4[ ������ � 02Dzh �������/ 
/@/./d/R/�/v/�/ �/�/�/�(���/?&? 8?J?�/n?\?~?�?�? �?�?�?�?O�?4O"O XOFOhOjO|O�O�O�O �O�O�O__._T_B_ x_f_�_�_�_�_�_�_ �_oo>o�/Voho�o �o�o(o�o�o�o�o (:Lp^�� ������ �6� $�Z�H�~�l������� ؏Ə��� ��0�2� D�z�h���To��ȟ� ��
���.��>�d�R� ������z�Я����� ��(�*�<�r�`��� ������޿̿��� 8�&�\�Jπ�nϐϒ� �������ϴ��(�F� X�j��ώ�|ߞ��߲� �������0��T�B� x�f���������� ����>�,�N�t�b� ���������������� :(^�v�� ��H���$ HZl:�~�� �����2/ /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?P?R? d?�?�?�?t�?�?O O*O�?NO<O^O�OrO �O�O�O�O�O�O__ 8_&_H_J_\_�_�_�_ �_�_�_�_�_o4o"o XoFo|ojo�o�o�o�o �o�o�o�?6Hf x���������v&��$TBC�SG_GRP 2�$�u� � �&� 
 ?�  Q�c�M��� q��������ˏ���*�1�&8�d,� �F�?&�	 H�CA�����b��CS�B��I�����V�>���d��n�Ќ�ԝB��g333��Blt�������AÐ�fcff:��.�C��z��l�?����G�w�R���A&��̧�����@��I��-� ��
�X�u�@�R������̻�����	V3�.00I�	mt	7���*� �%���ֶY��@ffj&� &�H�� N�� �O�  ����a� ϏϘ�*�J21��'8��Ϥ�CFG� )�uB� �E������d���#��#�I�W� �pW�}�hߡߌ��߰� �������
�C�.�g� R��v�������� 	���-��Q�<�u�`� r�����������I� cp"4��gRw ������	 -?�cN�r� �&������/ </*/`/N/�/r/�/�/ �/�/�/?�/&??J? 8?Z?\?n?�?�?�?�? �?�?O�? OFO4OjO XO�O�O`�O�OtO�O _�O0__T_B_x_f_ �_�_�_�_�_�_�_�_ ,ooPoboto�o@o�o �o�o�o�o�o�o( L:p^���� ���� �6�$�F� H�Z���~�����؏Ə ����2��OJ�\�n� ������������ �
�@�R�d�v�4��� ������ί����ү (�N�<�r�`������� ��ʿ̿޿��8�&� \�Jπ�nϐ϶Ϥ��� ������"��2�4�F� |�jߠߎ����߀���  �߼�B�0�f�T�� x����������� �>�,�b�P������� ��v�������: (^L�p��� �� �$H6 lZ|����� �/�/ /2/h/�� �/�/�/N/�/�/�/
? �/.??R?@?v?�?�? �?j?�?�?�?�?O*O <ONOOO�OrO�O�O �O�O�O�O _&__J_ 8_n_\_�_�_�_�_�_ �_�_o�_4o"oXoFo ho�o|o�o�o�o�o�o �/$6�/�oxf �������� ,�>���t�b����� ��Ώ��򏬏��&� (�:�p�^��������� ܟʟ�� �6�$�Z� H�~�l�������دƯ ��� ��D�2�T�z� h���Jȿڿ���� ��
�@�.�d�Rψ�v� �Ͼ����Ϡ����� �*�`�r߄ߖ�Pߺ� �����������&� \�J��n������ ������"��F�4�j� X�z�|����������� ��0B�Zl~ (������� ,Pbt�D�������   # &0/"��$TBJOP_�GRP 2*���  K?�&	H"O#,V,����� ��� =k%  ]Ȫ � �� �$� @ g"	 ߐCA��&��SC��_%g!�"wG��"k��/��+=�CS�?��?�&0~%0CR  B4�'�??J7�/�/?333�2Y&0}?�:;��Iv 2�1�0-1*20Ѽ6?�?20��7C�  D�!�,� B�L��OK:�Z�Bl  @pB@��� s33C�1 <�?gO  A�zG�2�jG�&)A)E�O�J;���|A?�ffY@U@�1C�Z0zjO�Oz@���U�O�$�fff0R)_;^;xCsQ?ٶ4)@�O �_tF�X_J\EU�_�VO:�t-�Q(B�*@ �Ooh�&-h$oZGLo 6oDoro�o~o8o�o�o �o�o3�oRl�Vd��V4�&`��q�%	V3.0=0m#mt7A@�s�*�l$!�'� �E��qE����E�]\E��HFP=F��{F*HfF@D��FW�3Fp?�F�MF����F�MF���F�şF���F�=F����G�G�.8�CW�RD3�l)D��E"���Ex�
E���E�,)F�dRFBFHFn�� F��F���MF�ɽF��,
GlG�g!G)�G=���GS5�Gi�Ĉ;��
;��o�|& : @�Xz&/��&�"�?�0�&=;-ES�TPARS  �(a E#HRw�AB�LE 1-V) I@�#R�7� � �R�R�R�'#!*R�	R�
R�R����!R�R�R�N��RDI��`!��@ԟ���
�r�Oz����������̯ޮ��Sx�^# <�����ÿտ �����/�A�S�e� wωϛϭϿ������� ;-w�{�_"��6��1� C�U���%�7�I�[�����NUM  V�`!� $ � ��m���_CFGG .���!@H �IMEBF_TT`}���^#��G�VE10�m�H�]�G�R 1=/�� 8�"� �� �A�   ������������ � 2�D�V�h�z������� ������/
e@ Rhv����� ��*<N` r������'/ //]/8/J/`/n/�/ �/�/�/r���_��t��@~�t�MI_CWHANS� ~� !3�DBGLVLS��~�s�$0ETHER_AD ?��w0�"��/�/�?�?l��$0ROUTq�!��!�4�?�<SN�MASKl8~�}1255.2E�s0OBO�TO�st�OOLOF/S_DI}��%V9�ORQCTRL C0���#��MT�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o�o&l�OIo8omoq�PE_DETAIJ8��JPGL_CON?FIG 6�����/cell�/$CID$/grp1qo�o�o/壀�?Zl~� ��C���� � 2��V�h�z������� ?�Q����
��.�@� Ϗd�v���������M� �����*�<�˟ݟ�r���������̯@�} a���&�8�J�\���^o��c��`���˿ݿ ���Z�7�I�[�m� ϑ� ϵ��������� �!߰�E�W�i�{ߍ� ��.����������� ��A�S�e�w���� <���������+��� O�a�s�������8��� ����'9��] o����F�� �#5�Yk}������`��User Vie�w �i}}1234567890� //,/>/P/X$� �cx/���2�U�/ �/�/�/??s/�/�3�/b?t?�?�?�?�??�?�.4Q?O(O:O@LO^OpO�?�O�.5O �O�O�O __$_�OE_�.6�O~_�_�_�_�_�_7_�_�.7m_2oDo�Vohozo�o�_�o�.8 !o�o�o
.@�o�agr l?Camera��o������ �ޢE �*�<�N��h�z���0�����I  �v�) ��$�6�H�Z�l�� ��������؟���� �2�Y��vP9ɟ~� ������Ưد����  �k�D�V�h�z����� E�W�I5����� � 2�D��h�zό�׿�� ��������
߱�W�ދ ��X�j�|ߎߠ߲�Y� ������E��0�B�T� f�x�߁ulY����� ����
����@�R�d� ��������������� W� iy�.@Rdv �/����� *<N��W��i� �������/ */</�`/r/�/�/�/�/as9F/�/?? 1?C?U?�f?�?�?D/ �?�?�?�?	OO-O�j	�u0�?hOzO�O�O �O�Oi?�O�O
_�?._ @_R_d_v_�_/OAO�p �{,_�_�_oo)o;o �O_oqo�o�_�o�o�o �o�o�_�u���oM _q���No�� �:�%�7�I�[�m� NEa����ˏݏ� ���7�I�[���� ������ǟٟ����ͻ p�%�7�I�[�m��&� ����ǯ�����!� 3�E�쟒�9�ܯ���� ��ǿٿ뿒��!�3� ~�W�i�{ύϟϱ�X� ����H����!�3�E� W���{ߍߟ����������������  ��L�^�p������������� ��   "�*�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/p`/r/�/�  
���(  �@�( 	 �/�/�/�/�/ ? ?6?$?F?H?Z?�?�~?�?�?�?�*2� �l�O/OAO��eO wO�O�O�O�O��O�O �O_TO1_C_U_g_y_ �_�O�_�_�__�_	o o-o?oQo�_uo�o�o �_�o�o�o�o^o poM_q�o��� ���6�%�7�~ [�m���������ُ ���D�!�3�E�W�i� {�ԏ��ß՟��� ��/�A�S���w��� ��⟿�ѯ����� `�=�O�a��������� ��Ϳ߿&�8��'�9� ��]�oρϓϥϷ��� ������F�#�5�G�Y� k�}��ϡ߳������ ����1�C�ߜ�y� �������������	� �b�?�Q�c������ ��������(�) p�M_q������0@ �������� ��#f�rh:\tpgl�\robots\�m10ia4_7l.xml�Xj |�������.��/1/C/U/g/ y/�/�/�/�/�/�/�/ /?-???Q?c?u?�? �?�?�?�?�?�?
?O )O;OMO_OqO�O�O�O �O�O�O�OO _%_7_ I_[_m__�_�_�_�_ �_�__�_!o3oEoWo io{o�o�o�o�o�o�o �_�o/ASew �������o� �+�=�O�a�s�����@����͏ߏ�I� �<<;  ?��4� �,�N�|�b������� ʟ�Ο���0��8� f�L�~���������������(�$TP�GL_OUTPU�T 9����� $�9�K� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ�����$�����2345678901��� �2� D�V�^����υߗߩ� ������w����'�9�K�]���}g���� ����o����1�C� U�g���u��������� ��}���-?Qc �������� �);M_q	 ������� %/7/I/[/m///�/ �/�/�/�/�/�/?3? E?W?i?{??%?�?�? �?�?�?O�?OAOSO eOwO�O!O�O�O�O�O��O_�O� $$Ӣ��OW=_o_a_ �_�_�_�_�_�_�_�_ #ooGo9oko]o�o�o �o�o�o�o�o�oC5g}��������}@��"��� ( 	  iW�E�{�i�����Ï ��ӏՏ���A�/� e�S���w�������� џ���+��;�=�O����s����Ƹ  <<\ޯ�)� ͯ�)��M�_���ʯ ����<���ؿ��Ŀ�  �~�$�V��BόϞ� x�����2ϼ�
ߤ��� @�R�,�v߈���p߾� ��j�������<�� ��r������� ���`�&�8���$�n� H�Z������������ ��"4Xj��R ��L���� |Tf ��v ��0B//�&/ P/*/</�/�/��/�/ h/�/??�/:?L?�/ 4?�??n?�?�?�?�?  O^?�?6OHO�?lO~O XO�O�OO$O�O�O�O _2___h_z_�O�_ �_J_�_�_�_�_o.o���)WGL1.�XML�cm�$T�POFF_LIM� Š�p����qfN_SVy` � �t�jP_M�ON :��ԍd�p�p2miST�RTCHK ;佥�f~tbVTCOMPAT�h*q�f�VWVAR <r�mMx�d � e�p�bua_�DEFPROG �%�i%MA�IN A_MES�A_IRVISI��`�rISPLA�Y�`�n�rINST�_MSK  �|� �zINUSE9R �tLCK)��{QUICKME�p�O��rSCREl����+rtps�c�t)������b��_桉STz�iRAC�E_CFG =��iMt�`	nt
�?��HNL 2!>�z���T{ zr@� R�d�v���������К��ITEM 2?�,� �%$12�34567890<�%�  =<�C�<U�]�  !c�k�wp'���ns�ѯ5� ���k������j�ů ��鯕���A�1�C�U� o�y�󿝿I�oρ�� ��	��-ϧ�Q���#� 5ߙ�A߽�����e߳� �����M���q߃�L� ��g��ߋ����%� w� �[���+�Q�c� ��o��������3��� {�;������G _����/�Se .�I�m�� �=�a/3/ ������k// �/�/�/]/?�/�/�/ ?�/u?�?�??�?5? G?Y?�?+O�?OOaO�? mO�?�?�OO�OCO_ _yO+_�O�Ox_�O�_ �O�_�_�_?_�_c_u_ �_o�_Wo}o�o�_�o o)o;o�o�oqo1C �oO�o�o��% ��[��Z���S�@��_�� 3 ے_� ����y
 Ï�Џ�~��UD1:\����q�R_GRP� 1A �� 	 @�pe�w�a�@��������ߟ͞�� ��ّ�>�)�b�M�?�  }���y��� ��ӯ������	�� Q�?�u�c���������Ϳ�	-���o��SCB 2B{� h�e�wωϛϭ���������e�UTORIAL C{���@�j�V_CON?FIG D{��������O�OUTP�UT E{�����������%� 7�I�[�m����� ���������%�7� I�[�m���������� ������!3EW i{������� �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/��/??'? 9?K?]?o?�?�?�?�? �?�/�?�?O#O5OGO YOkO}O�O�O�O�O�O �?�O__1_C_U_g_ y_�_�_�_�_�_�O�_ 	oo-o?oQocouo�o �o�o�o�o�_�o );M_q��� ���yߋ����-� ?�Q�c�u��������� Ϗ���o�)�;�M� _�q���������˟ݟ � ��%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ���
�� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� ��������������� 1CUgy�� �����	- ?Qcu��������/�x���$/6/ !/a/� �/�/�/�/�/�/�/? ?'?9?K?]?�?�? �?�?�?�?�?�?O#O 5OGOYOkO|?�O�O�O �O�O�O�O__1_C_ U_g_xO�_�_�_�_�_ �_�_	oo-o?oQoco t_�o�o�o�o�o�o�o );M_q�o �������� %�7�I�[�m�~���� ��Ǐُ����!�3� E�W�i�z�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�π�'�9�K�]�o�~���$TX_SCRE�EN 1F8%w  �}�~�@��������
���� m&��\�n߀ߒߤ߶� -�?������"�4�F� ��j��ߎ������� ��_����0�B�T�f� x������������� ��>��bt� ���3�W (:L^���� ����e/�6/�H/Z/l/~/�//�/��$UALRM_M_SG ?����� �/���/�/)?? M?@?q?d?v?�?�?�?�?�?�?O�%SEV7  �-EF�"ECFG H�Ż��  ��@�  AuA   ;Bȁ�
 O�� �ŨO�O�O�O�O__�&_8_J_\_jWQAGR�P 2I[K 0���	 �O�_� I�_BBL_NOT�E J[JT��l�������g@�RDEFPR�O� %�+ (%�MAIN�_2m% OVoAozoeo�o�o�o �o�o�o�o@�[�FKEYDATA� 1K�ɞPp 	jG���_������z,(�����(POINT � ]'�)�  OO�K T}@o�V�ND�IRECT��� ?CHOICEB����TOUCHUP ׏؏�'��K�2�o� ��h�����ɟ۟����#�5��Y��y���/frh/gu�i/whitehome.pngd�`����Ưدꯀ{�point���0��B�T�f���  |�look������ʿ�ܿ�}�indirec�(�:�L�^�p�>{�choic���@������������{�touchup�@0�B�T�f�x���{�arwrgϲ��� �����߁��)�;�M� _�q��������� �����%�7�I�[�m� �������������� ��3EWi{� ������ /ASew��r� �����/!/( E/W/i/{/�/�/./�/ �/�/�/??�//?S? e?w?�?�?�?<?�?�? �?OO+O�?OOaOsO �O�O�O8O�O�O�O_ _'_9_�O]_o_�_�_ �_�_F_�_�_�_o#o 5o�_Goko}o�o�o�o �oTo�o�o1C �ogy����P ��	��-�?�Q���u���������Ϗj�܋�u�܏�(� s��Q�c�r�,I����A�POINT � ]��9� OOK� Tß�}�ILT�ER۟�}�REE�ZE ���TOUCHUPG�H�s� ��~�����߯�د� ��9�K�2�o�V�����茿ɿ��whitehom�����%�7�I�X��poin�ߍϟϱ�����<`���look}���(�:�L�^���indirec|Ϙߪ���������choic���� �2�D�V�h��k�o�touchup�ߠ���������g�o�arwrg ��"�4�F�X�j�a��� ����������w� 0BTfx�� �����,> Pbt���� ��/�(/:/L/^/ p/�//�/�/�/�/�/  ?׿�/6?H?Z?l?~? �?�/�?�?�?�?�?O �?2ODOVOhOzO�O�O -O�O�O�O�O
__�O @_R_d_v_�_�_)_�_ �_�_�_oo*o�_No `oro�o�o�o7o�o�o �o&�oJ\n ����E��� �"�4��X�j�|��� ����A�֏����� 0�B�яf�x������� ��O������,�>��ټL������u�����q���ͯ��,������"�	� F�X�?�|�c������� ֿ������0��T� f�Mϊ�qϮϕ����� �����,�>�?b�t� �ߘߪ߼�˟����� �(�:�L���p��� �����Y��� ��$� 6�H���l�~������� ����g��� 2D V��z����� c�
.@Rd �������q //*/</N/`/��/ �/�/�/�/�/�//? &?8?J?\?n?�/�?�? �?�?�?�?{?O"O4O FOXOjO|OSߠO�O�O �O�O�OO_0_B_T_ f_x_�__�_�_�_�_ �_o�_,o>oPoboto �oo�o�o�o�o�o �o:L^p�� #���� ��� 6�H�Z�l�~�����1� Ə؏���� ���D� V�h�z�����-�ԟ ���
��.���R�d� v�������;�Я��� ��*���N�`�r���Ж������@���>�@������ 	��+�=��,)�n� !ߒ�y϶��ϯ����� �"�	�F�-�j�|�c� �߇����߽������ �B�T�;�x�_��� �O��������,�;� P�b�t���������K� ����(:��^ p����G��  $6H�l~ ����U��/  /2/D/�h/z/�/�/ �/�/�/c/�/
??.? @?R?�/v?�?�?�?�? �?_?�?OO*O<ONO `O�?�O�O�O�O�O�O mO__&_8_J_\_�O �_�_�_�_�_�_�_�� o"o4oFoXojoq_�o �o�o�o�o�o�o�o 0BTfx�� ������,�>� P�b�t��������Ώ ������(�:�L�^� p��������ʟܟ�  ����6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z����� -�¿Կ���
�ϫ� @�R�d�vψϚ�)Ͼπ��������*�`�,��`���U�g�y�Qߛ߭߇�,���ߑ����&�8� �\�C���y��� ���������4�F�-� j�Q���u��������� ���_BTfx �������� ,�Pbt�� �9���//(/ �L/^/p/�/�/�/�/ G/�/�/ ??$?6?�/ Z?l?~?�?�?�?C?�? �?�?O O2ODO�?hO zO�O�O�O�OQO�O�O 
__._@_�Od_v_�_ �_�_�_�___�_oo *o<oNo�_ro�o�o�o �o�o[o�o&8 J\3����� ��o��"�4�F�X� j��������ď֏� w���0�B�T�f��� ��������ҟ����� �,�>�P�b�t���� ����ί�򯁯�(� :�L�^�p�������� ʿܿ� Ϗ�$�6�H� Z�l�~�Ϣϴ����� ����ߝ�2�D�V�h� zߌ�߰��������� 
��.�@�R�d�v�ﴚ�qp���qp���������������,	N�r� Y������������� ��&J\C�g �������" 4X?|�m� ����/�0/B/ T/f/x/�/�/+/�/�/ �/�/??�/>?P?b? t?�?�?'?�?�?�?�? OO(O�?LO^OpO�O �O�O5O�O�O�O __ $_�OH_Z_l_~_�_�_ �_C_�_�_�_o o2o �_Vohozo�o�o�o?o �o�o�o
.@�o dv����M� ���*�<��`�r� ��������̏���� �&�8�J�Q�n����� ����ȟڟi����"� 4�F�X��|������� į֯e�����0�B� T�f�����������ҿ �s���,�>�P�b� �ϘϪϼ������� ���(�:�L�^�p��� �ߦ߸�������}�� $�6�H�Z�l�~��� ����������� �2� D�V�h�z�	��������������
�}�����5@GY1{�g,y �q���< #`rY�}�� ���/&//J/1/ n/U/�/�/�/�/�/�/ �/ݏ"?4?F?X?j?|? ���?�?�?�?�?�?O �?0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�_�_'_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o $�oHZl ~��1���� � ��D�V�h�z��� ����?�ԏ���
�� .���R�d�v������� ;�П�����*�<� ?`�r����������� ޯ���&�8�J�ٯ n���������ȿW�� ���"�4�F�տj�|� �Ϡϲ�����e���� �0�B�T���xߊߜ� ������a�����,� >�P�b��߆���� ����o���(�:�L� ^�������������� ��}�$6HZl ��������y  2DVhzQ��|�Q�����������,�/./�/R/9/v/ �/o/�/�/�/�/�/? �/*?<?#?`?G?�?�? }?�?�?�?�?OO�? 8OO\OnOM��O�O�O �O�O�O�_"_4_F_ X_j_|__�_�_�_�_ �_�_�_o0oBoTofo xoo�o�o�o�o�o�o �o,>Pbt� ������� (�:�L�^�p�����#� ��ʏ܏� ����6� H�Z�l�~������Ɵ ؟���� ���D�V� h�z�����-�¯ԯ� ��
����@�R�d�v� �������Oп���� �*�1�N�`�rτϖ� �Ϻ�I�������&� 8���\�n߀ߒߤ߶� E��������"�4�F� ��j�|������S� ������0�B���f� x�����������a��� ,>P��t� ����]� (:L^���� ���k //$/6/ H/Z/�~/�/�/�/�/h�/�/���+������?'?9=?[?m?G6,YO�?QO �?�?�?�?�?OO@O RO9OvO]O�O�O�O�O �O�O_�O*__N_5_ r_�_k_�_�_�_�_�� oo&o8oJo\ok/�o �o�o�o�o�o�o{o "4FXj�o�� ����w��0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� ����(�:�L�^�p� �������ʯܯ� � ��$�6�H�Z�l�~��� ���ƿؿ���ϝ� 2�D�V�h�zό�ϰ� ��������
���_@� R�d�v߈ߚߡϾ��� ������*��N�`� r����7������� ��&���J�\�n��� ������E������� "4��Xj|�� �A���0 B�fx���� O��//,/>/� b/t/�/�/�/�/�/]/ �/??(?:?L?�/p? �?�?�?�?�?Y?�? O�O$O6OHOZO�$U�I_INUSER  ���{A��  �[O_O_MENH�IST 1L{E�  (��@3�(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1�O__1_�C_�)�O�O527��@RRA_ESTEIRA�O�_�_�_��3'X_j^71�P_?PLACE0�_o�.o@o�9*�_jUed�it�BMAIN,22Lo�o�o�o�>�O�_955o-?Q�_�oq8
�����S_u�B422 �$�6�H�Z��o�p�3
o����ʏ܏�0���0�A����"�4�F�X�j� �������� şן�x���1�C� U�g�����������ӯ ������-�?�Q�c� u��������Ͽ�� ���)�;�M�_�qσ� ϧϹ��������� %�7�I�[�m�ߑߔ� ������������3� E�W�i�{������ ����������A�S� e�w�����*������� ����=Oas ���8��� '�0]o�� ������/#/ 5/�Y/k/}/�/�/�/ B/�/�/�/??1?C? �/g?y?�?�?�?�?P? �?�?	OO-O?O�?PO uO�O�O�O�O�O^O�O __)_;_M_8�O�_ �_�_�_�_�_�Ooo %o7oIo[o�_o�o�o �o�o�o�ozo!3 EWi�o���� ��v��/�A�S� e�w��������я� �����+�=�O�a�s��^[�$UI_PA�NEDATA 1�N������  	�}�  frh/cg�tp/flexd�ev.stm?_�width=0&�_height=�10ԐŐice=�TP&_line�s=3Ԑcolu�mns=4Ԑfo�nܐ4&_pag�e=doubŐ1���\V)  rim#�L�  ��c�u��� ������$�ϯ�گ� ��;�M�4�q�X����� ��˿�����%�\V�� � E�?  �b]���Dʟܝ2����2/�-�ual����_�� "�4�F�X�j�ώ�u� ���߫�������� B�)�f�M�������3�  I� ������*� <�N�`�����Ϩ��� ������i�&8 \C��y��� ���4Xj=��������� �� /S$/��H/Z/ l/~/�/�/	/�/�/�/ �/�/ ?2??V?=?z? a?�?�?�?�?�?�?
O }�@OROdOvO�O�O �?�O1/�O�O__*_ <_N_�Or_Y_�_}_�_ �_�_�_�_o&ooJo 1ono�ogo�oO)O�o �o�o"4�oXj �O������O ��0�B�)�f�M��� �����������ݏ� �>��o�o������� ��Ο��3��w(�:� L�^�p���韦����� ܯï ����6��Z� A�~���w�����ؿ� ]�o� �2�D�V�h�z� Ϳ�����������
� �.ߕ�R�9�v�]ߚ� �ߓ��߷������*��N�`�G����	��������������"�) ��G���6�s������� ����4������� K2oV���� ����#������$UI_POSTYPE  ��� 	 �/�UQUICKMEN  d�s�WREST�ORE 1O��  ��*defau�lt��  OU�BLE�PR�IM�mmen�upage,1422,10/d/v/�/��/=$editH"MAINQ/�/�/�/? ;%?4?F?X?j?|?! �?�??�?�?�?O "O4O�?XOjO|O�O�O CO�O�O�O�O_�?_ +_=_�Ox_�_�_�_�_ c_�_�_oo,o>o�_ boto�o�o�oU_�o�o �oMo(:L^ �����m� � �$�6��o�U�g�� ����Ə؏����� � 2�D�V�h��������xԟ�SCRE��?�u1�sc�u2�3��4�5�6�7r�8��TAT`�� ��MUScER�����ks����3��4��5��6ʨ�7��8��UND�O_CFG P�d����UPDX�����Non�e���_INFOW 1Q�<��0%��W���E���i� ��������տ��� :�L�/�pς�eϦύ�)�OFFSET Td@���{�� ����	��-�Z�Q�c� �߇ߙ��ϝ�������  ��)�V�M�_�q��������
���t���)�WORK U4�����A�S��Ͼ��UFRAM ����&�RTOL_�ABRT��$���E�NB����GRP �1V��Cz  A���+ =Oas������U������MSK � �<���N���%4��%��)��_'EVN�����>v�2W��
 h���UEV��!�td:\event_user\-F�C7���}�F�ցSP��sp�otweld�!C6����!�Z/�/:'�H/ ~/l/�/�/�/�/-?�/ Q?�/? ?�?D?�?h? z?�?O�?)O�?�?O qO`O�O@ORO�OvO�O _�O�O7_�O[__Z�]W+�2X����8V_�_�_ �_�_o �_,o>oobotoOo�o �o�o�o�o�o�o :L'p�]�����$VARS__CONFI�Y�˷ FP{���|C7CRG�\���>�{�t�D� BeH� pk�a�C�� ��}�?���C,&Qo=��ͩ�A ��MR2b����	}�	��@�%�1: SC130EF2 *����{�e����X� �5}������A@k�C�NF� w�Q�[� ��|����������T����\�ϟ �\� B���;� e�@�ǟ`�����S��� ��̯���ۯ�&�}� �\�G�Y���E���ȿ.�TCC�c
��h������pGF�p�gd��-�2�34567890�17�?��ׁ$��� 4�v�Nm�� ��϶��BW�����i�}�:�o=LA�څ�6��@�6�ͿZ���i�7����(��W���-�]�X� jĈߚߕϳϹ����� ����%�7�I�r�m� ߨ�ߵ��������� �8�3�E�W������ }��������������/�A�S�e�w��MO�DE��t �R?SLT e�|k�%"zς��;�1���d��`��SEGLEC��c��	�IA_WO�Pf� �� W,�		������G��P �����RTSYNCSE�� ��$�	#WINU�RL ?*ـ�;\/n/�/�/�/�/��uISIONTM�OU���A# ���%�gSۣ�S�ۥP�� F�R:\�#\DAT�A\�/ �� wMC6LOG?   UD16�EX@?\�' ?B@ ���2T1�  abriel?_Fariak?P5�?�?����� n6  ���GV<�2\� -��5��   ��Z�@�U058TRAIN�j?��*B{Rd_Cp|��D #`{2Х�'$�"��h#� (�kI�Mw��O�O�O �O�O1__U_C_]_g_�y_�_�_�_�(STA� i��@�o o2o�I8$>obo�%_GE��j#��~@ ��
�\��btgHOM�IN�kSۮ�B�`�2,,��CW���BveJMPER�R 2l#�
  ��I:��"�4F wj|�����`����&%S_g0�RE�m�^۴LE�Xdn�1-e�hoVMPHASE'  �e׃Bޱ�OFF _ENB�  �$VP2��$oSۯ��x�c C;�@ �a<;���?s33'D*AA��]� ��0ޱ�`r}�XC��܅���� ��[��6������6���]���>V�YD-۟E B��[�t\16���+FV���W��5d� ����,�>�'Es���`W�I�ǟ��� �� I�����9�k�ɯ;� ������ׯɿ3�տ�� ��C�8�g�Yϋ��ϯ� ��ϱϿ�����-�"� Q�c�u�jߙ�?��ϗ� �߻����u���M�B� T��u��߁����� ����7�,�[�m�� ]�k�}���������� !�E�����CUg ���!���� / !�-WQ��� ���c	//�)/?/M's�TD_F�ILTE�`s�k3 �x2�`����/ �/�/�/�/	??-??? Q?�6�/~?�?�?�?�?��?�?�?O OoiSH�IFTMENU [1t}<5�%5� ~O)�\O�O�O�O�O�O �O�O'_�O_6_o_F_�X_�_|_�_�_�_	�LIVE/SNA�P�Svsfli�v���_�z`I�ON ҀU
`bmenu&o+o�_�o�o�V"<E�uz��4IM�O�v���zq�W�AITDINEND  �ec��b�fsOKوOUTr�hSDyTIMdu��o|G�}#��{C�zb�z�xR�ELE��ڋxTM��{�d��c_AC�T`و��x_DA�TA wz���%�  EGA_BA�RRA_ESTE�IRA�o6Ex�RD�IS
`E��$X�VR�ax�n�$�ZABC_GRP� 1yz���� ,�2̏.MZD^��CSCH�`z����aP@�h@�IP�b{'���ş�ן�[�MPCF_�G 1|'���0 �r�8��� �}'�(�{p�s� 	(����  <l0 � ��
?� � 3�]9��5���ɓ���e3�[�����A  &Cj���D��a1w�?������{b?�7O��b�?�=.I�������2M\��������|2MPեǤ%Ϥ�ׯ7N 믙����o���w����� ˩�3����u�B� �˴2�۱�7�l �ĸǡ�	��1�?� i˟���ïբ0ۯQ���	��`~����_C_YLIND~!�� Р ,(  *.�?ݧ+�h�Oߌ�s� ������ ��(�	�x�-��&�c� �߇�������j�P� ���)��~�_�q���� �2�'��� � &����������&h��I��cA����SPHERE 2�������� ��A�T/A��e ������ /N`=/�a/H/Z/��/��/�/�/��ZZ� ��f