��   ��A��*SYST�EM*��V9.3�044 1/9�/2020 A� 
  ����DRYRUN_T�  4 $�'ENB  �$NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��SAW_� G �%$INIT�	RESUME_�TYPENDIS�T_DIFFA $ORN41� d �=R0�&J_�  4 $:(F3IDX���_ICI  ��MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_SIZc���� ��. h $USE_FLC 3!p�:&iF*SIMA�7#QC#QBn'SC�AN�AX�+IN��*I��_COUN�rRO( ��!_TMR_VA�g#h>�ia �'�` ����1�+W[AR�$�H�!��#N3CH�P�E�$O�!PR�'I�oq7iOq ��OoATH-� P $ENA#BL+�0B�T�$$C�LASS  ����A��5��5��0VERS�G�  fAIRTU� O@'/ �@E5���"����-@{FA@A�E��%A�O���O�Ob����QEI2\K�*_<_N_`_r_�_ �_�_�_�_�_�_oo�&o8oJo�O*W?<"Hg@ ���j�@�o�o�i�� � �2\I  4%Xo��}A�A�o ;_qP������@�A���� 8��)�n�M�A@�c$"P+ �k�K-@��ń�AЄX�A@A-@�N ��
��.�@�R�d�v� ��������П���F�A 偍A��(�:�L�^� p���������ʯܯ��DxL	|W� 2���h�O�a�s� ��������Ϳ߿�� �'��A�Z�l�~ϐ� �ϴ���������� � 2�=�V�h�zߌߞ߰� ��������
��.�@� K�d�v������� ������*�<�G�Y� r��������������� &8JU�n� ������� "4FXc|�� �����//0/ B/T/_q�/�/�/�/ �/�/�/??,?>?P? b?ah�4�0���?�p