��   �;�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����DCSS_CPC�_T 4 $�COMMENT �$ENAB�LE  $M�ODJGRP_N�UMKL\  $UFRM\~] _VTX M ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�? �ELAY_T�IMJSPEED�_CTRLKOV�R_LIM? p JD� L��0�UTOO�i��O���&S. � 18J\TC�u
 !���\�� jY0  �� �CHG_S{IZ�$AP!��E�DIS�]$!�C_+{#s%O#)J�p 	]$Jd#�  �&s"�"{#�)�$�'��_SEEXPA�N#N�iGST�AT/ DF�P_BASE �$0K$4!,� .6_V7>H73h}J- � }܏\AXS\UP�LW�7���9a7r �< w? �?�?��?�?�//�	7ELEM/ �T �&B.2NO0�G]@%CNHA�DF#~� $DATA)qhe0  P�J�@ 2 
:&P5 �� 1�U*n   _VS iSZbRj0jR(�VyT�(�R%S{TROBOT�X�SARo�U~�V$CUR_���RjSETU4"	� �bAISP_M�GN�INP_ASSe#�PB!� `C iH�77`e�.fXc1��CONFIG_wCHK`E_PO* �}dSHRST�gM�^#/eOTHERRBT�j_G]�R�d�Tv �ku�chT1r
0R HLH�d� 0 � lt<Ne'AV�RFYhH^t�5�1ȕ ��W�_A$�R��UPH/ (G%Q�Q�Q�3wBOX/ 8�@F!�F!�G �r�{�zTUIRi@ � ,�F�pE}R%@2 $�po L�_SF�� "�ZN/ � IF(@�p��Z	_�0�_�0wu0  @�Q7yv	
��~  �$$CL`  �������Q��Q��VER�SION���  0��IRTUAL���'� 2 �Q  G�p���&@)>�m�����������������Ғd<��Cz  0�� ��A���l��������� Ɵۯ���� �2�D� F�h�}�����ԯſ�� ���
��.�@�R�d� fϋϚ�����п���� ���*�<�N�	�rχ� �Ϩ�b��Ͼ����� &�8�^�\�n߃��� ����������"�4� F�X�m�|������ �������0�B�h� Vx����������� �,>Pbw �������/ /(:L�`/��/ ����/�??$/ 6/H/Z/l/�?�/�?�/ �/�?�/�?O#O2?D? V?h?jO�?�O�?�?�? �O�O__.O@OROdO vO�O�_�_�O�O�_�O 	oo�_<_N_`_r_-o �_�o�_�_�o�_�o )8oJo\o�o�o�o� 2�o�o��o�%�4 FXj|������ ������!�3�B�T� f���z�������ҏ� ����/�>�P�b�t� ��������Ο����� �+�=�L�^�p���� ����ʯܯ���'� 9�H�Z�l�~����ϴ� ��ؿ����#�5�G� V�h�zόώ߰����� ������1�C�R�d� v߈ߚ߬߮������� 	��-�?���`�r�� ��Q����������� ;M\�n������� ���V����"7 IXj|���� ����/E/W/ fx���/��/� �/?,/A?S?b/t/ �/�/�/�?�/�?�/? O(?=OOOaOp?�?�? :O�O�?�O�? OO'_ 6OK_]_lO~O�O�O�O �_�O�_�O_#o2_Go Yokoz_�_�_�_�o�_ �o�_
o@o1 Ug vo�o�o�o�o�o�� -�<Q�c��� ���u����� Ώ8�*�_�q��������ʏȏڋ�$DCS�S_CSC 2����Q  P����:�܉d
�k�.���R��� v�ׯ����Я1��� U��y�<���`���ӿ �������޿?��c� u�8ϙ�\Ͻπ��Ϥ� �����;���_�"߃� Fߧ�j߷��ߠ���� %���I��m�0����f��������GR�P 2�� ����	ҟS�>�w�b� �������������� =(aL�p� �����  K6oZ�~�� ����/5/ /Y/ D/}/h/�/�/�/�/�/ �/?�/
?C?.?g?R? �?�?�?z?�?�?�?�? O-OOQO<OuO�O�O dO�O�O�O�O_�O_ ;_&___q_�_N_�_�_ �_�_�_�_�_%ooIo���_GSTAT �2��%��<� ����2?�S��?̓?�� 5�Y׵�T׵鼠�`���S��¶���C��MD#���8`<�e��߸?t�䁴��0.����` ��a>�`4��Z�/1�Cv������e>�	y�m��Q>xN�=��̾m|u�x�\�iB�U]�Ρ�C~ y�=�>龢W!�?q�޿t���`´�g{>��w�f�f�����C����V�C�S y������:?WnU`pmdpghp��?u�&>o��>>"뫴`�C��XD�j y���z?K}�?	���p�o��J�"�5� Ϳ�`�`�a��o �o�ov��<�N���0� z���f���Љ�i�a -i��+k y �.��&� H�v�\�~�������� ȟڟ��*���Z�l��� x���|���د���.� �B��J�0�B�d��� x���ȿ��������� �F�H��Ϻ�tϾ���Ϫ�����͵����?�6<�R��b5��t��j߷��P4�޿��5@�K�C�"D)���m�<rE�?����b���1�~���bqмm��a@���C���m�M�q�YR?���� gʿ��ٿYe������ó`C��� y��Q>���� ?r�;��q�<rDN�����eњ�r��p������������C��ް�ڌ�-���>��:�e�� �p���pK&����@�MC��ߑDB�� y<p�]�?�)<��MJ���<pK�9��/5��}�I�0�O�F�(�:�L� ���������� ���� V�h��Pϒ�dϪ��� ��������F, ^|bt��j�� 8��<N(r� z�������� �,//4/b/H/Z/|/ �/�/�/�/�/�"?T ?X?j?D?�?�?z?�� ��P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��O�?�?�?�?t_ �_|?�_�_�_�_�_o ��/.o ?FodoJo\o ~o�o�o�o�o�o�o �o2`?���_ ����� �od J�xB�d���x���ȏ ��Џ������F�,� N�|�b�(�������� ���*�<��4_F_�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ ~�`�r�����"�� .�X�2�DώϠ�:��� �Ϝ��� ������H� .�P�~�dߖߴߚ߬� ���ߢ�,�>�p�*�t� ��`���� ���� �� �.��6�d�J�l� �������������� ����Z��F��| ���п⿈����� ��Я�����*�<� N�`�r�������/�  ��/�/��/�/ �/�/*?<?��$f?8 ~?�?�?�?�?�?�?�? O O2OPO6OHOjO�O >�O�O?�O_"_�O F_X_N?�O�_�Oz_�_ �_�_�_ o�_o6oo .oPo~odo�o�o�o`_ �o(_�o,>bt Nl/~/$6HZl ~������� / /2/D/����� VH�Z�Pf���j�|� Ɵ؟r_�o��o�8� �0�R���f������� ί�ү��4��od� v���b���������� �8��L��8�f�L� nϜςϤ��ϸ����� � �"�P�6�����Ŀ ~����ߴ������� �������,� >�P�b�t��������� Ώ��R�4�F�X����� ����,bt �\ߞp߶��� �$R8j� n���v� //D �H/Z/4/~/�/�� �/��/�/?�/
?8? ?@?n?T?f?�?�?�? �?�?�?�/.O`/OdO vOPO�O�O�O����\� n����������� ���"�4�F�X�j�|� �_�O�O�O�O�o�o�O �o�o�o�o�o�/�? :ORpVh�� �����$�
�� >�l�O�����o��� ��Џ�,�"p�V��� N�p�������ԟ��ܟ 
���$�R�8�Z��� n�4�ʯ���� ����6�H�V��$DCS�S_JPC 2�@�Q (G D1������� ��P��ۿ������ ��Y�(�g�Lϡ�p� �ϔ��ϸ����1� � �g�6�H�Z߯�~��� ���������?�� � u�D�V�h������ ���)���M��.�p� ��d�v��������� ��7[*N� r�����!� /i8�\�� �����//�/ "/w/F/�/j/�/�/�/ �/?�/�/=???0? �?T?�?x?�?�?�?�? O�?�?8O]O,O>O�O bOtO�O�O�O�O�O#_ �OG__k_:_L_�_p_��_�_�_�_�_��h�S
q�u�L�_Uooyo��dDo�oho�o�o�o �o�o1�oUy @Rd����� ��?��c�*���N� ��r�����󏺏̏ޏ ��M��q�8���\��� ��ݟ���ȟ%���� �Y��F���j�ǯ�� 믲��֯3���W�� e�B���f�x������� ����A��e�,ω� Pϭ�t��ϘϪϼ�� +���O��s�:ߗ�^� �߂��ߦ������� K��$�6�H��l��� ��������5���Y�  �}�D�V�h������� ������C
g. �R�v���� ���Qu<� `����/�&d�MODEL 2�3kx��
 �<�c (  �z(�/g/y/�/ �/�/�/�/�/�/D?? -?z?Q?c?u?�?�?�? �?�?�?.OOO)O;O MO_O�_�OY/�O�O_ �O�O<__%_7_�_[_ m_�_�_�_�_�_�_�_ 8oo!onoEoWo�o{o �o�o�o�o�o�O�O�O �o|�oew�� ����0���+� =�O�a�������䏻� ͏ߏ���b�9�K� ��3Es����m�۟ ����#�p�G�Y��� }�������ůׯ$��� �Z�1�C�U�g�y��� ؿ����ϩ������ h��Q�cϰχϙ��� ���������d�;� Mߚ�q߃��ߧ߹��� ����N�%�7��� 1�C�q��Y�����&� ���\�3�E�W�i�{� ������������ /A�ew�� ��������� =O�s���� ���/P/'/9/�/ ]/o/�/�/�/�/?�/ �/:??#?5?�?/ ]?o?�?�?�?O�?�? HOO1OCO�OgOyO�O �O�O�O�O�O�OD__ -_z_Q_c_�_�_�_�_ �?
o�?�_�_Ro)o;o �o_oqo�o�o�o�o �o�o<%7I[ m������� ��!��_��oI�[� ȏ������Տ���� �/�|�S�e������� ����џ�0���f� =�O�a�s�����m��� ����ѯ>��'�t�K� ]�o��������ɿۿ (����#�p�G�YϦ� }Ϗ��ϳ�����$��� �����5�Gߴ�/� �߯�������2�	�� h�?�Q�c�u����� ���������)�;� M���q�����k�}߫� ��*��%7I[ ������� �\3E�i{ ����/��F/ ����!/3/�//�/�/ �/�/�/?�/?T?+? =?O?�?s?�?�?�?�? O�?�?OPO'O9O�O ]OoO�OW/i/{/�O�O �O�O_^_5_G_�_k_ }_�_�_�_�_o�_�_ Hoo1oCoUogoyo�o �o�o�o�o�o�o�OV �O1u��� �
�����)�;� ��_�q���������ˏ ݏ�<��%�r�I�[��m����$DCSS�_PSTAT ����ӑ�Q    l�� � (��+��O���t�  r�Ԑ�������������ӕ௎�կ�Ĕ�SETUP 	NәBȖ����� 8�R�ͬs�b����������T1SC 2
4+�����Cz�������صCP R�D�DLj�|� >�ϲ��ϓ������ ��0�B�T�#�xߊ�Y� �����ߡ������� >�P�b�1����y� �������(���L� ^�p�?����������� ������$6Zl ~��Vϫ�D�� �);Mq� �d����// �7/I/[/*//�/�/ r/�/�/�/�/?!?�/ ?W?i?8?�?�?�?�? �?�?�?�?O/OAOO eOwOFO�O�O�O��O �O_�O+_=_O__s_ �_�_f_�_�_�_�_o o�_9oKo]o,o�o�o �oto�o�o�o�o# �oGYk:��� ������1� � �g�y�H��������� ���	��O-�?�Q�؏ u�����h���ϟ��� ���;�M�_�.��� ����v�˯ݯ����� %���I�[�m�<����� ����ٿ���̿!�3� �W�i�{�Jϟϱ��� ���������/�A�S� "�w߉��j߿��ߠ� ������=�O�a�0� ����x������� �'���K�]�o�>��� ��������������# 5Yk}L�� �����1C gy�Z߯�� Z�	//�?/Q/c/ 2/�/�/h/z/�/�/�/ ??)?�/M?_?q?@? �?�?�?�?�?�?�?O %O7OO[OmOONO�O �O�O�O�O�O�O�O3_ E__i_{_�_\_�_�_ �_��_oo�_AoSo eo4o�o�ojo�o�o�o �o+�oOas B��x���� �'�9��]�o���P� ����ɏ�����Ώ#� 5�G��k�}���^��� şן�������_C� U�ܟ6�����l���ӯ 寴�	��-���Q�c� u�D�����z�Ͽ�� ¿�)�;�
�_�qσ� RϧϹψϚ������ %�7�I��m�ߑ�`� �����ߨ������3��E�W�&��$DCS�S_TCPMAP  ������Q @ U.�.�.�.ક�.�.�.��.�	.�
.�.��.�.�.�/� � .�.�.��.�.�.�.�T.�.�.�.�.�U.�.�.� .�U!.�".�#.�$.�U%.�&.�'.�(.�U).�*.�+.�,.�U-.�..�/.�0.�U1.�2.�3.�4.�U5.�6.�7.�8.�U9.�:.�;.�<.�U=.�>.�?.�@u�UIRO 2����������� ����,>Pb t�������-���-��Qc u������� //)/;/M/_/q/�/ �/2�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O�/3O �/WOiO{O�O�O�O�O �O�O�O__/_A_S_�e_w_�_�_&O�_q�U�IZN 2��	 ����� oo$o *��_Rodovo9o�o�o �o�o�o�o�o*< Nr��Y�� ����&�8��\� n�=�������ȏ��� ���ߏ4�F�X��|� ����o�ğ֟蟫�� �0���T�f�x�;�M� �����������_x�UFRM R�����81�^�p�/� ������ʿܿ�� �� �6�H�#�l�~�YϢ� �Ϗ��������� �2� I�V�h�ߌߞ�y��� �߯���
���.�@�� d�v�Q������� �����*�A�N�`��� ����q��������� ��8J%n�[ ������" 9�FX�|�i� ����/�0/B/ /f/x/S/�/�/�/�/ �/�/??1(?P?b? =?�?�?s?�?�?�?�? O�?(O:OO^OpOKO �O�O�O�O�O�O __ )?;?H_Z_�O~_�_k_ �_�_�_�_�_�_ o2o oVohoCo�o�oyo�o �o�o�o
3_@R �ov�c���� ���*��;�`�r� M�������̏ޏ��� �+8�J��n���[� ������ǟ���ٟ"� 4��X�j�E�����{� į֯������