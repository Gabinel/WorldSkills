��   v��A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����UI_CONFI�G_T  x� L$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY73��ODE�
4CF�OCA �5CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%��!BA�!j ��!BqG�#�!hINSR�$IO}7PM��X_PKT?�$IHELP� M�E�#BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�<STY.f2$Iv!_Gv!�k FKE�FHT�ML�_NAM��#DIMC4:1]ABRIGH83s oDJ7�CH92%!FEL0T__DEVICg1&�USTO_@ o t @AR$@'PIDD�BC�D*7PAG� ?hA�B��ISCREuEF����GN�@$FwLAG�@��&��1  h 	$�PWD_ACCES� MA�8��hS:1�%)$LAB=E� $Tz j�HP�3�R�	4SU�SRVI 1  < `�R*�R�n�QPRI�m� �t1�PTRIP�"m��$$CLASP ����a��R2��R `\ SI�	g�  0�aIRTs1	o`�'2 L1�L1���R	 ,��?���a1`��b�d~a���� � �`y�o��
 ��a��o�o1CU  �oz�����c �
��.�@�R��v� ��������Џ�q�� �*�<�N�`���� ����̟ޟm���&� 8�J�\�n��������� ȯگ�{��"�4�F� X�j���������Ŀֿ����`TPTX�����/�`� sȄ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ��� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F�X���|��������������a�f�b�� ($p�-����T�?�x���a�a��c���c����l��c�g���aR�ah�ah��at2�h�	f�����������a���`  ����f ep)��h#h�F�bc� Xc�B 1)hR_ \ _�� REG �VED]���w�holemod.�htm�	sing}l	doub �trip8?browsQ� ����u����//@/���d/ev.sl�/3� 1�,	t�/_�/ ;/i/??/?�/S?e?pw?�?�?�?� � �?�?OO%O7OIO[OmOO�E @�?�O�O �O�O�O_�F�	�?�? ;_M___q_�_�_�_�_ �_�_�_oo%o7oIo [omooM'�o�o�o�o �o�o+=Oa s������� ��?>�P�b�t����� ����Ώ���O��� ��L�^�_'_����� ��ş�����6�1� C�U�~�y�����Ư�� ӯ�o���-�?�Q� c�u���������Ͽ� ���)�;�M�_�-� �ϬϾ��������� *�<�7�`�r�A�Sߨ� ��q���i�����!� J�E�W�i����� ��������"��/��� O�I�w����������� ����+=Oa s������� ,>Pbt�� �߼���//�� ���^/Y/k/}/�/�/ �/�/�/�/�/?6?1? C?U?~?y?�?Y��?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__�R_d_v_�_ �_�_�_�_�_�_�o�*o�_o`oro�j�$�UI_TOPME?NU 1K`�a�R 
�d�a*Q)*de�fault5_]�*level0{ * [	 �o��0�o'rtp�io[23]�8?tpst[1[x)�w9�o	�=h5�8E01_l.p�ng��6mencu5�y�p�13�z���z	�4���q��]���������̏ޏ )Rr���+�=�O�a�~��prim=��page,1422,1h�����şן ����1�C�U�g����|�class,5p�����ɯۯ�����13��*�<��N�`�r���|�53�������ҿ�����|�8��1�C�U�g�y� ���ϯ���������"Y�`�a�o/��m!ηq0�Y��avtyl}T�fqmf[0nl�	>��c[164[w�Ճ59[x�qG�y��tC	8�|�29��o�%� 1���{��m��!��� ��0�B���f�x���`������o���80��'9K~���2 P�����\�� '9K�������������1���/$/6/H/Z/U�~|�ainedi'���/�/�/�/�/P�c�onfig=si�ngle&|�wintp���/$?6?H?�Z?	�ߐ??ٷ�gl[57�ٳq��?�;$gp�08�ݲ07I�?hF��F2JO[6�:��?)O�O�x �� �4s�x�O���$� �`�o�H_Z_l_~_�_ �_Q��_�_�_�_o o �_DoVohozo�o�o�oz�!;�$doub5�o��13��&du�al�i38��,4�o&�o9�o�n�o �a8���Ao�����&�8��%3L=}!��o�b8@����� ����z���(�:���+:T��i48,2�o��b{����ʟ  {?�;�M�sc���;����s�� �}���e�u0��X��@�F7L���@`�O��2�h�z�6e�u7�����ｿϿ�0��̏�27��G� Y�k�}Ϗ��0�s�Ϡ�������!�1 �M�_�q߃ߕ���� ���������7�I� [�m���������@�����!�����6(��]�o��������$��746�����)�C��ߟT�	TPTX[209�<AwA2IHJ���Bw1H��]H�����02��A#��[T�tv`��O�L#_�0� \��5S[�tre�eview3v�3���~�381,26 M/_/q/0�/�/�/ �/�/�/~/?%?7?I? [?m?�o/(��o5%����?�?�?�A�?\1~��?8"2��eOwO�? �?(}�LEK��O�O_ �O��8@�ONOa_s_�_��6_d�E_�_�_�_ oV�#_���_�Sooo �o�oB�o�o��oA �oq+=Oa s��o����� ��(�9���Q�x��� ������ҏ?���� ,�>�P�ߏt������� ��Ο]�����(�:� L�^�ퟂ�������ʯ ܯk� ��$�6�H�Z� �l�������ƿؿ� y�� �2�D�V�h��� �Ϟϰ������ϕo�o ��o@ߧE�c�u߇� �߽߬�����O���� )�<�M�_�q���W� ��������&�8��� \�n���������E��� ����"4��Xj |����S�� 0B�fx� ���O��// ,/>/P/�t/�/�/�/ �/�/]/�/??(?:? L?��߂?1ߦ?�� �?�?�?�?O$O5OGO �?SO}O�O�O�O�O�O �O�O��2_D_V_h_z_ �_�_�/�_�_�_�_
o o�_@oRodovo�o�o )o�o�o�o�o* �oN`r���7 �����&��J� \�n���������E�ڏ ����"�4�ÏX�j� |�������a?s?蟗? �sO_/�A�S�e�w� ������������� �,�=�O�a�#_���� ��ο��=��(�:� L�^�pς�Ϧϸ��� ���� ߏ�$�6�H�Z� l�~�ߐߴ������� ����2�D�V�h�z� ������������
� ���@�R�d�v����� )���������ƚ�Ԕ*defau�lt%��*level8�ٯw����? tpsOt[1]�	�y��tpio[23���u���J�\menu7__l.png_|13��5�{�y4�u6���/ /'/9/K/]/���/�/ �/�/�/�/j/�/?#?�5?G?Y?k?�"pr�im=|page,74,1p?�?�?��?�?�?�"�6cl?ass,13�?*O@<ONO`OrOOB5xO@�O�O�O�O�O�#L �O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]ooo��o`�$UI_U�SERVIEW �1֑֑R 
���o��o�o[m�o' 9K] ���� �l���#�5��o B�T�f������ŏ׏ 鏌���1�C�U�g� 
���������ӟ~��� ��v�?�Q�c�u��� *�����ϯ�󯖯� )�;�M�_�
��~��� ���ݿ���%�ȿ I�[�m�ϑ�4ϵ��� �����Ϩ�
��.ߠ� i�{ߍߟ߱�T����� ����/���S�e�w� ���Fߨ����>�� �+�=�O���s����� ����^�����' ����FX��|�� ����#5G Y�}����p ���h1/C/U/g/ y//�/�/�/�/�/�/ �/?-???Q?c?/p? �?�??�?�?�?OO �?;OMO_OqO�O&O�O �O�O�O�O�?�O_ _ �OD_m__�_�_�_X_ �_�_�_o!o�_EoWo io{o�o0h