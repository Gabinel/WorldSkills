��   2�A��*SYST�EM*��V9.3�044 1/9�/2020 A� 
  ����PASSNAME�_T   0 �$+ $~'WORD  ? �LEVEL  �$TI- OUT�T  &F/�� $SETU�PJPROGRA�MJINSTAL�LJY  $�CURR_O�UwSER�NUM��STSTOP_T�PCHG V L�OG_P NT��N�  6 COUNT_DOWN��$ENB_PC�MPWD� $D�V_� IN� s$C� CRE��MA RM9� T9DIAG9(��LVCHK F�ULLM/�YX=T�CNTD��MENU�AUT�O+�FG_DS]P�RLS�U�BURYBAN�v!/8&ENC/�  CR�YPTE ~�  �$$CL(   ���K!���	��	@ V� I�ONH( � 0�\!IRT�UA� J/�$DC�S_COD?�|��O%�  W�'q_� �/�(S  �*%�� � �&�A9�1�"�!	 $R!�� =,?B? P?f?t?�?�?�?�?�? �?�?OO(O>OLObO\��3SUP� :a�dOvO3F�O��O�O��  �\Q��&_ ��� V�[t&�+�j��T�O~_ ��<W:_��t �V�_�GLUGH 1�)_ t �) oo'o9oKo]ooo�o �o�o�o�o�o�'�_	 -?Qcu�� �����o��)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ���/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� �������� ��'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� ��
��1�C�U�g�y� ��������������	 �-?Qcu�� ������%