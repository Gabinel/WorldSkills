��   ��A��*SYST�EM*��V9.3�044 1/9�/2020 A� 
  ����DRYRUN_T�  4 $�'ENB  �$NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��SAW_� G �%$INIT�	RESUME_�TYPENDIS�T_DIFFA $ORN41� d �=R��&J_�  4 $:(F3IDX���_ICIfMIX�_BG-y
_�NAMc MOD�c_USd�IFoY_TI� ��MKR-  �$LINc  { "_SIZc�� �. h �$USE_FL�C 3!�:&iF*S�IMA7#QC#QB�n'SCAN�AX֋+IN�*I��_C7OUNrRO( ���!_TMR_VA�g#h>� ia �'` �����1�+WAR�$ҵH�!�#N3CH��PE�$O�!PER�'Ioq7iOq�fOoATH-� P $ENA#BL+�0B�Tf�$$CLA�SS  ����A��5��5�0V�ERS�G�  0�AIRTU� O@'/ �@E5���"����-@{FA@A�E��%A�O���O�Ob����QEI2\K �O;_M___q_ �_�_�_�_�_�_�_o�o%o7oIo�O)W?y"Hg@ �� �j@�o�o�i�� �� 2\I  #4%Xo��}A�A �o;_qP������@�A��� �8��)�n�M�A@�c�$"+ �k�K-@��ń�AЄXV�@A-@ �N��
��.�@�R�d� v���������П���F �A偍A��(�:�L� ^�p���������ʯܯ��DxL�W� 2�l�O�a� s���������Ϳ߿� ��'��A�Z�l�~� �Ϣϴ����������  �2�=�V�h�zߌߞ� ����������
��.� @�K�d�v����� ��������*�<�G� Y�r������������� ��&8JU�n �������� "4FXc|� ������// 0/B/T/_q�/�/�/ �/�/�/�/??,?>? P?b?ah�4�0���?�p