��   ?Q�A��*SYST�EM*��V9.3�044 1/9�/2020 A�   ����MN_MCR_T�ABLE   �� $MACR�O_NAME %$PROG@�EPT_INDE�X  $OP�EN_IDaAS�SIGN_TYP�D  qk$M�ON_NO}PR?EV_SUBy a �$USER_WgORK���_L� �MS�*RTN �  &SOP�_T  � {$�EMGO�}�RESET��MOT|�HOL�l��12�S�TAR PDI8�G9GAGBGC��TPDS�RE�L�&U� �� �EST��^�SFSP�C����C�C�NB���S)*$8*$3�%)4%)5%)6%)7�%)S�PNSTR�z�"D�  �$$�CLr   �S���!����� VERSION�(�  0���!IRTUAL��/�!;LDUIM�T  ��� ����4MAXDR)I� ��5
4.�1 �%� � d%Op�en hand 91����% ?�? �"  13�0?Closeo?�?��?	O�9�7Rel�ax�?�?GOmO�9�6j82oOPO�OtO�3�?�O�O&_�O�6 @+O__�_;_�4�F �_�_�_�_�[�3��(@ �_6o�_Zo	oo�o?o �o�ouo�o�o�o �o �oVS�;M� q����.��R� ����7���[�m��� �ߏ�ǏُN���r� !�3�m���i�ޟ���� �ß8�J���3���/� ��S�e�گ��ׯ��� ѯF���j��+����� ��ֿ����ϻ�0�߿ �+�x�cϜ�K�]��� ���ϥϷ���>���b� �#ߘ�G߼���}߷� ��(�����^��[� ��C�U���y����� $�6�!�Z�	����?� ��c�u������� �� ��Vz);u� q����@R ;�7�[m� ��/��N/�r/ !/3/�/�/�/�/�/�/ ?�/8?�/�/3?�?k? �?S?e?�?�?�?�?�? �?FO�?jOO+O�OOO �O�O�O�O_�O0_�O �Of__c_�_K_]_�_ �_�_�_�_,o>o)obo o#o�oGo�oko}o�o �o(�o�o^� 1C}�y��� $��H�Z�	�C���?� ��c�u�ꏙ�� �Ϗ �V��z�)�;��� ��柕����˟@�� �;���s���[�m�� �����ǯ�N���r� !�3���W�̿޿��ǿ �ÿ8����n��k� ��S�e��ω��ϭϿ� 4�F�1�j��+ߠ�O� ��s߅߿����0��� ��f���9�K���� ������,���P�b� �K���G���k�}��� ����(����^� 1C������ $�H�	C�{ �cu��/�� 	/V//z/)/;/�/_/ �/�/�/�/?�/@?�/ ?v?%?s?�?[?m?�? �?O�?�?<ONO9OrO !O3O�OWO�O{O�O�O _�O8_�O�On__�_ A_S_�_�_�_�_�_�_ 4o�_XojooSo�oOo �oso�o�o�o�o0�o �of�9K�� ����,��P�� �K�������k�}�� ���ŏ׏�^���� 1�C���g�ܟ�ן $�ӟH���	�~�-�{� ��c�u�ꯙ����ϯ D�V�A�z�)�;���_� Կ����Ͽ��@�� �v�%Ϛ�I�[ϕ��� ��ߵ���<���`�r��!�[�
Send �Events�S��SENDEVNT��Q���� %=	��Data�߶�ODATA��ڝ���%��SysVayr;��SYSVw���ڳO�%Get<�x�GET+������%Requ�est Menu����REQMEN	U?��۶�]ߞ�Y� ��}�+�����.�� d�7I�m ����*�N� ����i{� �/��/\/G/�/ //A/�/e/�/�/�/�/ "?�/F?�/?|?+?�? �?a?�?�?�?O�?�? BO�??OxO'O9O�O]O �O�O�O___>_�O �Ot_#_�_G_Y_�_�_ �_o�_�_:o�_^oo oYo�oUo�oyo�o  �o$6�ol� ?Q�u���� 2��V��������� q��������ˏݏ �d�O���7�I���m� ⟑���ݟ*�ٟN��� ���3�����i���� ���ïկJ���G��� /�A���e�ڿ����� "��F����|�+Ϡ� O�aϛ�����߻��� B���f��'�a߮�]���߁ߓ��$MAC�RO_MAXX�~���������SOPENB�L ��� 2��ݐѐ�_���"�?PDIMSK�2�3<�w�SU����TPDSBEX S K��U)�2� ����-�