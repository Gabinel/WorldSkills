��  	��A��*SYST�EM*��V9.3�044 1/9�/2020 A�  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���A�IO_CNV�� l� RAC�L�O�MOD_TY]P@FIR�HA�L�>#IN_OU��FAC� gIN�TERCEPfB�I�IZ@!LR�M_RECO"�  � ALM�"EkNB���&ON�!� MDG/ 0� $DEBUG�1A�"d�$3AOp� ."��!_IF�� � 
$ENABL@C#� P �dC#U5K�!MAЧB �"�
� OG��f 0CURR_tD1P $Q3LIN@tS1I4$C$AUSO�d�APPINFwOEQ/ ��L A ?1�5/� H �79E�QUIP 2n�0NAM� ��2�_OVR�$V�ERSI� �ST~�0COUPLE, �  $�!PP�V1CES0�!H1��!�PR0�2	 �� $SOFT��T_IDBTO�TAL_EQ� �Q1]@NO`BU SP?I_INDE]uE�XBSCREENu_�4BSIG�0�O%KW@PK_�FI0	$T�HKY�GPANE�hD � DUMM�Y1d�D�!U4� Q!RG1R�
 � $TIT1d ��� 7Td7T� �7TP7T55V65V7*5V85V95W05W>W@�A7URWQ7UfW1pW1zW1�W1�W 6P~!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$�Nb_OPT�2p��(CELLSETUP  `�0�HO�0 PRZ1%�{cMACRO�bR'EPR�hD0D+t@���b{�eHM M�N�B
1�UTO�B U�0� 9DEVIC&4STI�0�� P@�13��`BQdf"VA�L�#ISP_UN9I�#p_DOv7IyFR_F�@K%D1�3�;A�c�C_W�A?t�a�zOFF_�@N�DEL�xL�F0q�A�qr?q�p�C?�`�A�E1�C#�s�ATB�t��d�MO� �sE � [M�s���2�REV�BIL�F��1XI� %�R o � OD}`~j�$NO`�M�+��b�x�/��"u�� ����!X��@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQCw ��a_EDu >� � C2�e�`S�p�4%$l ��t$OP�@QB�qy�_OK���0, P_C� y��dh�U ^�`LACI�!�a��� FqCOMM� �0$D��ϑ�@�pX��OR BIG�ALLOW� �(KD2�2�@VA�R5�d!�AB e`BL8[@S � ,KJq�M�H`S�pZ@M_Ox]z���CFd7 X�0GR@�z�M�NFLI�<��;@UIRE�84<�"� SWIT=$/0k_No`S�"CFd0�M� �#PEED��!�%`����p3`J3tV�&$E��..p`L��ELBOF� �m��m��p/0��CP�� F��B����1��r@1J�1E_y_T>!@Բ�`��g���G�� �0WARN�Mxp�d�%`�V`N�ST� COR-�rFLTR�TR�AT T�`� $ACCqM�� R�r$ORI�.&ӧ�RT�SFg C�HGV0I�p�T(��PA�I{�T�!���� � p�#@a���HDR�B
��2�BJ; �C��U3�4�5�6�7�8�9>���x@ޮ2 @� TR�Q��$%f��ր��F��_U���ѡ�Oc <� ����Ȩx3�2��LLECM�}-�MULTIV4�"$��A
2q�CHI�LD>�
1��z@T_�1b  4� S�TY2�b4�=@�)�24����@�� A|9$��T�A�I`��E��eTO���E��EXT���ᗑ�B��22�0>��@��1b.'��}!9�A�K�  �"K� /%�a��R���?s!>�O�!M��;A�֗�M8�� 	�  =�I�" L�0[�� �R�pA��$JOB`B�����`���IGI�# dӀ����R��-'r��A�ҧ��_M���b$ tӀFL�6�BNG�A��TBA� ϑ�!��
/1�@À�0���R0�P/pX ����%�|���Bq@W�
2JW�_)RH�CZJZ�_*zJ?�D/5C�	��ӧ��@��Rd&A������ȯ�qGӨ�g@NHANC��$LG/��a2qӐ� ـ�@��A�p� ���aR���>$x��?#DB��?#RA�c?#AZ�t@�(.�����`FCT����_F࠳`�SM��!I�+lA�% ` �` ���$/�/�@���[�a��M�0�\��`��أHK��A�Es@͐�!�"W��Nz� SbXYZW�`D�"����6��C�����'  . I�I��2�(p�STD�_C�t�1Q��US�TڒU�)#�0U�[�%?IO1��� _Up�q�* \��=�#AORzs8Bp�;�]��`O6  RSY�G�0�q^EUp��H`�G�� ��]�DBPX�WORK�+���$SKP_�pAqf�au@�TR�p , �=�`����Z m�OD3��a _�C"�;b�C� �GPL :c�a�tőS�D�W�3Bb����P�6�P )DB�!�Y-�B APR��
I�8Ja3��. /�u�\���� �LuY/�_ȔS��0�_����PC�1�_�TEN9EG�]� 2�_�S�VPRE.��R3H� $C��.$L8c/$uSނz IkgINE�WA_D1%�ROyp�������`�q�c7 t@�fPA��~�RETURN�b.��MMR"U��I�;CRg`EWM@�/SIGNZ�A ����e� 0$P�'�1$P� m�	2p�p'tm�+pD�@ �'�bdNa)r�GO_AW ��h@ؑB1�@CSd��(�CYI�4���`1Pw�qu��t2�z2�v�N�}��E}sDE�VIs` 5 P7 $��RB���I�wPk��I_B�Y���"�T7Q�tH�NDG�Q6 H�4��1�w��$DSBLC��o��vg@��4I�qL��7O�f@�]���FB���FE�ra8�ׂ�t}s���8�> i�T1?���MC�S���fD �ւ[2H� W��EE���%F�p���t����9 T�p<��x�NK_N:���j��U��L�wHA�v	Z' ~�2���P~r��q7: �=MD	Ln���9�ጂٱh�����!e����J ��~�+����,�N�D����3��ՒG!aq�SLAd�7;  ��INP��"�����X}q_ �4<�06`�C� NU��  jD�Lק��SH!�
7=M��q���ܢ�Ӣ���g���>P +$ٰ�٢���^��^�Y�FI B\��Ă��'A	r'AWl�NTV��r]�V~�X�SKI�#�T���a�ۺ�T1J�3:3_�P�SAF�N���_SV�EOXCLU��N@�%DV@Ll @�Y����S�HI_V
0\2P�PLYPRo�HI�M�T�n�_MLX�>�pVRFY_�ClM��IOC�UC!_� ����O�qţLS�0v�FT4Q������@P�E$t�t��A��CNFt��6եu��pm�4ACH�D�o������AF&C CPlV�TQTP8?�� �� ?`�@�TA�@�0L@ r��N��]� @����T��T! S����t<e@{RA DO�� �w2���!$n��_1�#�H!�̔��΀K��B�2��M/ARGI�$�����A ��_SGNE�C;
$�`�a ^aR0��3��@ B��|B��ANNUN�P@?���uCN@�`�%0����� ���BEuFc@I�RD @Q�1F���4OT�`�s�FT�HR,Q��CQ0�M��NI|RE���r��AW���DAY=CLOAD�t;T|�<S�5}�EFF_AX�I��F`1QO3O���Eq��@_RT+RQE�G����0+RQj�Evp ��|�F�0f�R0 ��t �AMP�E><� H 0�``œ^�`Ds�DU�`����BCAr� �I?�`N ErID?LE_PWRI\4V!n0V�wV_[ |྅ �DIAG�5J�� 1$V�`SE�3TQl�e��0Pl�^E_��j��VE� �0SW�H�q(� �b|�G�n�OHxPPLHk�IRAl�B�@ �[��a�bk��w3��O � ��v�|�I��0 �pRQDWf�MS-�%AX{<6j�LIFE�@�&�MQy�NH!Q%��$F#C����CB0��mpN$�Y @�aFL�Al���OV0]&H�E��l�SUPPO$�@u�y��@_�$�冀!_X83�$gq�'Z�*W�*B1�'T�#`�fk2XZáj�Y2D8ECY`T@�`N����f� �C�k����ICTA�K `�pCACH�ӫ�3з���I��bNӰUFFI� \��@���;T��<S6CQ.�MS�W�5L 8	�KE�YIMAG�cTM La��*Ax�&E���B��OCVIER-aM; ��BGL����y�?� 	��П4�N�:�ST�!�BP�D,P�D��D<��@EMAI䐔ax��M�s�FAUL|RAObB�c�� spUʰ�MA"`T'`E�P<' $S�S[ � ;ITw�BUF�7y��7�tN[�LSUB1T�Cx�o�R�tRSAV|U>R'c2�\�WT���P�T�*`�Sn�_1PbU���YOQT�bK��P��M��d���WAX��2���X1P��S_GH#
?$�DYN_���Q <Q�D��0��U�M�� T�eF�`|�\�DI�ҏEDT_Pɰ:�R$��b�GRQM�&��Jq��a���׀��Fs� oS (�SVqp�B��4�_�.��a��T� �@���Bn�SC_R]1IK>B'r��$t��R"A#u�HN�aDSP:FrP�lyIM|Sas�qz��aB� U>w� <1%sM�@�IP��s��0`tT!Hb0ЃTr��T`assHS�cCsBSCʴq0� V�����S�{_D��CONVE�AG���b0^v1PFH�y�dCs�`&a?ASC8���sMERg��a�FBCMPg��`E�T[� UBFU&� DU%P�D�:1�2�CDWy�p�P�CGM�[@NO6�:�V� ��� ���P���C"�����w��A��|`��WH *�LƠ�Cc�W����Y� 賂��р�q�|�P��A��7}�8}��9}�H ���1��1���1��1��1ʚ1�ך1�1�2��2T����2��2��2��U2ʚ2ך2�2�3��3��3����3���3��3ʚ3ך3��3�4��QEX	T[�X[b�H``t&�``z�k`˷$���F{DR�YTP�V��RK"	��K"R�EM*F��]"OV�M:s/�A8�TRO�V8�DT�PX�MX�g�IN8ɉ W��INDv�["
�ȕ`K ^`G1a�a��@Q%79Da�RIV��u"�]"GEAR:qIO.K(�[$N�`����,(�F@� \#Z_MsCM<0K! �F� 9UT���Z ,�TQO? b�y@t�.G?t�E |�p.�>Q����[ �5Pa� RI�E���UP2_ \ �@=STD	p<T�T���������a>RB;ACUb] T��>R
�d)�j%C�E��0��IFI��0��i�{��4�PTT��FLU=I�D^ �?0gHPUR�gQ�"�r�aP�4P+ I�$��]Sd�?x��J�`sCO�P�SVRT��>N�x$SHO* ��CASS��Qw%�pٴBG_%��3��࣓��FOR�C�B��o�DATAZ��_�BFU_�1�b�b�2�en�b0��` �|K`NAV	`)������$�S�Bu#?$VISI���2SC	dSE������V��O�$&�B�K�� ��$PO���I��FM�R2��a  ��	��`#��@&�8�O� (�_��9��+IT_^�ۄ�)M�����DGC{LF�DGDY�LD����5Y&��Q$RY�M됇CbN@{	? T�FS�P�D�c P��W�cK �$EX_WnW1P%`]��"X3�5�s�G+�d �K`ָ�SWeUO�DE�BUG��-�GRt��;@U�BKU���O1R� _ P�O_ )�����M���LOOc>!SM E�R�a��u _E� e >@�G_�TERM`%fi'��ORI�ae gi&�`SM_�`>Re !hi%V�(ii%3�UP\Bj� -����e��w#� f���G�*ELTOr�A�bF�FIG�2��a_���@�$�$g$wUFR�b$�01R0օ� OT_7F��TA�p q3NST��`PAT�q�0�2P'THJ�ԀE�@�c3ART�P'58�Q�B�aREL�:�aSHFT�r�a�1�8E_��R��у�& � 	$�'@i�
����sN@bSHI�0�Uy�= �QAYLO�p� Oaq�����1����pERV��XA��H�� m7�`�2%�P�E3�P��RC���ASYM�a��aWJ07����AE�ӷ1�I��ׁUT@�`Oa�5�F�5P�sXu@J�7FOR�`M &P�GRO!k]��`5&�0L0���HOL ;l �s2T�����OC1!E��$OP��qn����$�����$��PR�^��aOU��3e���R�5e�X�1 �eo$PWR��IMe�BR_�S�4�� �3��aUD���`�Q�dm���$H�e!�`AWDDR˶HR!G�2��a�a�aQ�R��[�n H��S����%��e`3��e���e��SEl��L�HS�MNu�o���Pªq��0OL�s߰`ڵ�I ACRO��&1��ND_C�s��Afd�K�ROUP��R_�В� �Q1|�=�s ���y%��y-��x���y���y>�=A��Ҁ�AVED�w-��u�`<(qp $_��P�_D�� ��'rPR�M_��HTT�P_�H[�q (�ÀOBJ��b �$˶LE~3�P��\�r � ���ྰ%_��TE#ԂS�PIC��KRLPiHITGCOU�!��L�� �PԂ������PR��P�SSB�{�JQUE?RY_FLAvs�@_WEBSOC��G�HW�#1��s�`}<PINCPU(���O���g�����d�t��O��IO�LN�t 8��R���$SL!$INPUT_U!$`��Pw�֐SSL.���u����2�.��C��B�IO^a�F_AS=v��$L+ਇ+�A ��bb41�����Z@�HYʷ����#qe�U;OP:w `v�ϡ�˶�¡�������"`P IC`���� �	�H��IP_ME��v�x Xv�IP�`(�R�C_N�p�d���R0ʳp�ױQrSP �z��C��BG(� ��M��Av�y lv@CTiApB��AL TI�`3UfP_ ۵�0PSڶBU_ ID� 
�L �� `�a�����0�z)����ϴ�N�N�_ O��IRCA�_CNf� { ��Ɖ-�CYpEA��������IC����tpR�=QDAYy_
��NTVA������!��5����SCAj@��CL�
����
���v�|5�VĬ2,b�l�N_�PCV�n�
���w�})�T��S�р���
��e���T� 2| $� �v��~��֣�ذLABp1��_ ��UNIX�9�ӑ ITY裪�D�ea�R� ��<)����R_URL���$A;qEN ���ts`vsTeqT_U���J��X�M�!$���E�ᒐR祪�"� A�,���JH���#FLy��= 
����
�UJR|U� ���F�6G��K7��=D>�$J7�s��J8*�7���3�E��7��&�8\�)�AP�HIQ4�y�D�kJ7J8R��L�_KE'�  ��K͐LMX� 7� <U�XRi������WATCH_V�AZqu@AំFIE�L`��cyn���:�� � u1VbwPC�TX�j�����LGE��� �!��LG_SIZ�΄�[8Zm�ZFDeIYp1!gX b ZW �S`�8� m��� �b ��A�:0_i0_CMc3#�*'FQ1KW rd(V(Bb�po pm�p� |I�o�1 pb pW RyS��0  (C�SLN�R�۠�DE6E3����c��i���PL#�DAU"%EAq�͐�T8"�. GH�R��y�BO�O�a�� C��F�ITV�l$A0��sRE���(SCRX�����D&�ǒ�qMARGI4�Sp�,�����T�"�y�S��x�Wp�$y�$��JGM7�MNCHt�y�FNĤ�6K@7r�>9UF�L87@L8FWDL8H]L�9STPL:VL8�"�L8s L8RS�9HOPh;��C9D�3R��}P�'IUh�`4�'��5$ ��S2G09�pPOWG�:�%�3,64��vN9EX��TUI>5I� �ӌ�����C3�C<0'�,�o:��&��@�!NaqvcANAy��Q�AI]�gt7���DCS���cRS�c*RROXXOdWS�ÂRroXS{X�(IGNp �
Ђ=10 ��[TDE-V�7LL��Y"*��C �	 8�Tr$@f/蛒����3A�a�	 W�萦�Oq�s�S1Je2Je3�Ja��BSPC � �ƋG`-T��%���Q�T�r@�&E�fST��R9 YBr�a /�$E�fC�k��g��f	v9�CB� L����� ��u�xs뀀��g�q�jt��!�#_ ���ʐv�#Ӽ� �s �MC��� ���CLDP|᠜�TRQLI ����y�tFL���rQ���s5�D���w~�LD8�u�t�uORG���1��RESERV���M���M�Œ�t��� � 	�u�5�tF�uSV��p��	1������RCLMC���M�_�ωА��_C��MDBGh�I�����$DEBUG�MAS������U��$T8P��EF�d��pFRQҤ� �� K	HRS_KRU4�bq��A���$EFREQ6u!y$0YOVER�Ђk��f�PU1EFI�%Gq�� �7�9
Y�z�� \�����E�$U�`��?���
�PSI`��	���CA ��ʲ�σU|Y�%�?( 	���MISC�� d���aRQ��	��TB� � ���A���AX��𑧪�EXGCESg�9d�M�
H�9�u���}qd��SC�` � H�х�_�����������pKE��+�� �&�B_, FLIC�BtB� QUIRE CMOt�O��얩quLdpMD� �p�{!��5b���$L��MND!��I�����L �D;
$I�NAUT�!
$RSM�ȧPN�b�Cx���PSTLH�w� 4U�LOC�f�RI"��eEX��A�NG.R.���ODA]��q��� �RMF0����icr�@pmu���$�SUPiuv��FX��IGG! � ���cs� �#cs
Fct��ޒ�b5� �`E��`T�5�tC��g&�TI��C`נ� �M���� t�M	D���)��XP��ԁ���H��.���DIAa��Ӻ�W�!��0af�*��D@#)֡O�㥀n��� �CUp �V	���.���O�!_��� �{`�c��L���� |�P|�h�0� ��P{�KEB��e-$B��o�=p�ND2ւ����2_{TXltXTRAXS4������LO: �1���}�L���C�.�&�[�RR2>h��� -�!�A�� d$CA�LI���GFQj�2�F`RINbn�<$Rx�SW0ۄ���wABC��D_J��{�q��_J3��
���1SP, �q�P�����3��H�9pq�B#J�3n���O�Q�IM耯�CSKP �zb7?SbJ+ᯂ�Qb�y����_cAZ��/�EL�Q<.ցOCMP�ð��� RTE�� �11�0 ���1��@: ZSMG�0��v��JG�pSCLʠ��SPH_�P���f��q�u�RTEIR��n�Pk�_EP
�q�`A� �c���sDI�Q23Ud�DF  ���LWn�VEL�qINxr�@�_BLXP.���Y/�J��'$ � �IN���]�C�9%�".�8!6p_T� �F%a"����^$��k)�~pDH�ʠ��\�9`$V0w��_�A$=��l~�&A$��S��h��H �$B�EL� m��_ACCE� 	8�0OIRC_�q�@��NT��c$PSʠ�rL���M4�s 9 .7��GP/6��9�7D$3�73S2T�͡_Ga��"�0�1��8�1_M�G}�DD�1�~�FW�p��3�5$32�8�DEKPPABN6[7ROgEE�2Ka BO�p�Ka��1�?$USE_v�S]P��CTRTY4@�� �� <qYNg�A �@�FR �ѢAM:�N��=R�0O�v1�DINC(��B�4���GY.��ENC�L��.��K12��H0IN�bI0S28U��ONT�%NT23_�~�fSCLO�~�|P��Iذ ~��V�~�$��hpU�#�CQ MVMOSI��1<�[�1����PERCH  �S��� �W���SlщR��l�@���E�0�0PAS2EeL�DP7�ONU�8�Z�f�VTRK�RqAY"�?c��aS2�e��c�����BP�MOM�B���C�H�}�C�j��c�3gBT�DU�X �2S_BCKLSH_CS2Fu:��V ���C-�esRoz�A�CLALMJT@��`� �uCHKe ����GLRTYpн�8Tȗ�5���_�ùT_U	M3��vC3��1Z�n��LMT��_LG��%���0�E*�K�=� )�@5F�@8 9�Nb��&)hPC�Q)hHТ��5�uCMC���0�7CN_��N���;SF�!iV�B��.W����S2/�ĈCAT�~SH�Å��4 V�q�/q/V�T1��0P�A�t�B_P�u�c_ f Z�f�Pe�cݔ�u�JG���ѓ�OG|އ�TORQU~@ �S�i @e��R� @B�_Wu�d�!a�P�#`��#`�Ih�Iv�I�#F��S�:��I�0VC00��֢�1ܮ�0��JRaKܬ!��<�DBX�Mt�<�M�_DL�!_bGRVg�`��#`��#A�H_%�?��0���COS��� ��LN#���ߥŴ� ��=@������꼰�<�Z���VA�MYǱ:ȧ���|��[�THET0�UNK23�#���#Ȱ[CB��CB�#Cz�AS�ѯ����#��Ɗ�SB�#��GT	SkZAC����x&���$DU�p@hg6�j��E�%Q%aY_��x�NEhs1AK�t�� y�A}��կ׍�����LPH����^U��Sߥ��� �������!��(Ʀ�EV��V�غ ��V��UV��V
�V�V&�V4�VB�H������P��d�����H
�H�UH&�H4�HB�O�ܥO��Os���O��O���O
�O�O&�O
4�O(�F�Ҫ�	����SPBALA�NCE_J�6LE6��H_}�SP>!۶�^�^��PFUL�Cb�q���K*1=�UTO_�p�u�T1T2�	
22N �q2VP�M�a� i�(Z23	qTu`O�1>Q�INSEG2�Q�REV�PGQDI�F�ep)1�U�1��`OBK�qj�w�2,�VP�qI�LCHgWAR4B�BAB��~u$MECH���J��A��vAX�aP�o���׫"� � 
p�?�10UROB�P�CRS2#%Ղ�@�C�1_ɒT � �x $WEIGH�@�`$��\#���I�A�PIFvA�0LAG�B��S�B:�B7BIL�%OD�`�P&s"ST0s"P:�pBt � N�C!L �P �
P2�Aɑ  2y��Tx&DEBU�#�L|0�"5�MMY�9C59N��$4�`3$D|1 a$0ې�l� > DO_::0AK!� <_ �&�� �q�A��B�"� N�JS�8_�P�@��"O��p �� %"�T7P?Q�TL4�F0TICK�#�TE1N0%�3=p�0N�P� u3�PR\p�A��5���5U0PROMP��CE�� $I�R"��A�p8BX`wBMCAIF��A�BQE_� COCX�a�@RU�7COD�#FU�@�&ID_�P�E82B> �G_SUFF�� ��#�AXA�2D�O�7/�5� �6GR �#��DC�D��E���E-��DU4� �_ Hn_FI�!9GS7ORD�! R 2�36s�HR�AN0$�ZDT�E=!� X5��4 *WL_N�A�1�0�R�5DEF_I�X�RF�T�5�"��6�$�6�S�5�UFISm�#�m1|��40c�3�T6�44􁆂�"�D� ?rfd�#D�O|@ l2LOCKE����C�?OG2a�B�@UM�E�R�D�S�D�U�D >b�B�c�E�S�Dd�B �&2v2a�C�ʑ�E�R��E�S�C9wwu�H�0P@} d�0,a��F0W�h��u�c480�T�E�qY4� >�!LOMB_�r�w�0s"VIS��IT�Ys"AۑO�#A_�FRI��~SI,a�n�R�07��07�)3�#s"W�W�Q���%�_���AEAS {#�B��|�x`WB8��45�55�6|#OR�MULA_I����G�W� h �
>75COEFF�_O�1&)��1��Gdo�{#S� 52CA� �:?L3�!GRm� ?� � $�`�v2X�0TM�g���e��2�c��3ERIT��d�T� �  �L�L�Dp`S��_SVLkd��$�v� �.����� � ��SE;TU,cMEAG@�@�Πt �!HRL � �3 (�  0��@l��l��aw��R�0$�a�a}d]�d��B��Ay`Gax`��[�:�k@REC[Qq���QSK_A y��� P_!1_USER�����*���VEL����-��!��IzPB�MT�1CFG��� � �0]O�NO#REJ �0l���[�?� 4 e���"�XYZ<SB� �3�0��_ERR�K!� U ѐ�1�@�c�Ȱ�!�>�B0B?UFINDX���P�� MORy�� H_ CUȱ�1��dA�yQ?�I>Q$ +�a����� \��G{�� � $�SI�h��@2	�V�Ov�q�- OBJE<| w�ADJUF2y�F��AY�����D�ǃOUKP����AMR=�T��-���X2DIR����Xf�1  DYNt�0�-�	T� ��R��0� �ҿ�OPWOR�� ��,B0SYSsBU����SOPo�H��z�Uy�XP�`K���PA�q����V��OP�@U����}�"1��IMAGb۱_ �п"IM.����IN������RGOVRD"ё�	���P����  >gplcC��L�`BŰ?l�P�MC_E�P�1N"��Mr�1212R��"�SL| ��� �^R OVSL=S�rGDEX\a`��2�:�_"���P#���@P������2�C �P>���#�_ZE�Rl���:���� �@��:��O�@RIy��
[�g@e���s��P�PL���  �$FREEY�E�U�~�Z��L�����T�� ATUSk�,1C_T�����B������p�Vc1���P��� Dc1�к���LQ����MQ��ۡL�XE��x�5IbP�W�` ��UP��H`&aPX;@��4y3����PGY�}�g�$SUB����q���JMPW�AIT~ ���LO�W���1wē CVF_A�0��R�Z���CC �R$��28I�GNR_PL��D�BTB� P*a�B�W@.t�U�0-I�G��!@I�TNL�N,�RBѡb�N<!@��PEED~ ��HADOW� ��t����E������PS�PD��� L_ A`�нP���	#UNq Ȫ �RP (�LY�wPa����PH_�PK���b�RETGRIE��x���2��R!D@FI��� �x��V �$ 2�d��DBGLV<LO�GSIZz�baKT�U���$D��_[TXV�EM�Cڡ�)�� �-R�#�r��CHECKz����L�J��ϰq)�L��.��NPA�`TJ"�����)1P����
�A�R�"�BC =Sa��O8�@����ATTS�u�䡳&� w�^a�3-#U1X^�4�PL�@Z��� $d��qSWI�TCH�h�W��A�S��f�3LLB���� $B�A�Dvc��BAM�i��6I��(@J5ȸ�N�UB6[F
A_KGNOWK3qB"�U��#AD+Hc� D��I?PAYLOAq�9pB�C_���GrѼGZ�C�LqAj��PLCL=_6� !4��BPOA?�T7�VFYACӐ�Jp��D�I�H!RՐ�G�TB��6��J(�zQ_J�A �B�AND����T�B�Q�����PL~@AL_ ��0� =�TAe��pC��D:�CE���J3�P�V�� T�PDCK�^�)b��COM�_AgLPH�ScBE<�߁�_�\�X�x\�� � ���OD�_1�J2�DDM�A�R<�h�e�f�cQ�TWIA4�i5�i6��MOM(��c�c�c�c4�cV�B� AD�cv��cv�cPUBP�R �d<u�c<u�b}"�1����� L$PI $��pc��G�y��I*�yI�{I�{I�s�`@�A���v��v�J��b��a��HIG �3���0���5 �0�f�?�5N�5�SAMPD Ƣ�0�p���;@�S �� с6���1���� �� �`���`1�K�P��`�d�P�H��IN1� �P��8�T�/��:�z�xQ�z���GAMM&��S��$GET������D^d>�
$N�PIBR��I��$HI��_���1��E=��A�9�*�LW�W�N�9�{�*��Zb���QCdCH�K0�j�ݠnI_ ��M�JļRoh�Q ���sJ�-v��S {�$�X 1�N�}I�RCH_D�$RN���^�L�E��i�p�Zh8�ž�MSWFL/Mn�PSCR�75��� ��3�"Ķ�6��`���ع�紙��0SV��P'�������GRO�g�S_SaA=AH�=ńNO^`Ci�_d=��no�O �O�x�ʚ��p�B�u���cDO�A��!� ں�*�t�:�Z1f�;��7����CFMmu� 7� �YL�snQ ��� ���"��<s�	�����nQ૰�<3M_Wl��� ��\p��(�o�MC��P���Q�����hpM.�pr� ���!��$�WM��ANGL�!�AM�6dK�=dK�DdK��TT7�N�k@��3�#�PXC O�Ec�QZ��hp	nt�[ ���OM��� ϑϣϵ����`� c��Z0es^a_�2� | a�J��i���c���c�J��j�����jA� O ,x��� ��@{�P�1�PMO�N_QU�� �{ 860QCOU�n�QTHxHO��nB HYS�0ESPBFB UE- 3�f0O�4�  c P�^��RUN_TO��rI�O��� P�@x��INDE�#�_PGRA���0��2>��NE_NO���ITf��o INF�O��a"�����vH�OI� (*�SLEQ!�*�*��Q OS��l4�{ 460ENABy�>� PTION�3�p�r��^GCF�!� @60J�Q���R�d!���erPEDIT�ԓ �� ��KAQ"�� �E(�NU'(A�UTY�%COPY�AQ�2,�qe�M�Nx< @+��PRUTm� C"N�OU�2�$G��$RGAkDJ��u2X_��AIX����&���&W�(�P�(~��&9�� 
�N^�P_CYCy�e1/RGNSc�{�s��LGO£�NYQ__FREQSrW@��X1�4�L�@�2P0p�!�c@�"�CRE���MàIF�q�NA���%�4_Gf�S�TATU~�f��M'AIL��|CIq�=�LAST�1a*4EwLEMg� ��Q>rFEASIt;� ւΰ��B"�F�AF����I� ��O2�E� u�vBAB��PE� =�VA�FzQ�I��bTqU[��R��S~�FRMS_TRpC �Qc��C��Z�
��1�Dc I�,2ns؆��	MB 2�  `���N�3V�R2WR*����шR^W�wj�DO�U�^�N�,2PR�`�h�1GRID���BARS!�T�YuZ�Op��+ |_�4!� �R�TO��d� � 9����POR�c\~vbSRV�0)"dfDI[�T�`;aNd�pXg
�Xg4Vi��Xg�6Vi7Vi8:av�F�ʒg�z $VACLU�C0�3D1AC�a>d�� !pf����S�1-ȆAN�/��c�0R�]11AT�OTAL����=sP�WE3I�QStREG#ENQzfr��X�H�0]5	v( TR�CS��Qq_S3��wfp�V �!��r��BE�3�P�G0B�( sV_H��PDA(��p�S_�Ya���i6S��AR�(�2� �"IG�_SE�3�pb�5_� �tC_�V$CMYPl��DEp�G�
��IšZ~�X�
���Fm�HANC.'� p Qr�2����INT9`cq�F<���MASK�3�@OVRMP �PD���1-��W�QaХT��l�_RF�{�V�PSSLGP�g�9� j5��,�;pDpS���4���U��.�}�T9E���`���`k�ⵥJ^�Y�y3IL_�Mx4�s��p��TQ@( ���@����V.��C<�P_ �R�F�M�]�V1\�V1j�2�y�2j�3y�3j�4y�4j���p۲�������ܲIN�VIAB8�6�#��*�2&�U22�3&�32�4&�!42��6���SJ�  ��T $MC�_FK `� �LP>�J�х1pMj�Iу��zS ��1����KEEP_HNA�DD��!鴓@�C��0	��Q����
�O!�v ���p
�և.
�REM!�	�CqP�RF�]�b�U�4e	��HPWD  ��SBM���PCOLLAB*�p��/q�2IT/0��Q"{NO1�FCALp�܎���� , �FL|v�A$SYN����M��Ck��RpU_P_DLY��z�DELA9�Dq�2Y� AD(�3��Q�SKIPO�� �4`� O��NT����c�P_� ��׾ �� cp���q�ٞ��o`�� |`�ډ`�ږ`�ڣ`����`��9�!�J2RT0  �lX�@TR3 H��1AH� �H����.�RDCq���+ � R�R, 5���R�1��E��5TR�GE�_C��RFL�G"���W�5TSsPC�1UM_H��2TH2N}Q��;� 1� ��;��Q02 �� D� ˈ��@2_PC3W�S���1Y0_L10_Cw2x��-��� � $ \� U@��V7������0��VU\��`��� rd��C *�T�7��DZ Gs�.RUVL1[�1h���v10]�_DS��������PK 11�� lڰ����q��AT?��$�Q[7�� ���K 5T���H7OME� ��c2h�n����(�&0`3h���0!3E *�c4h�hz�����5h���	/P/-/?/W6h�b/@t/�/�/�/�/�7h��/�/??'?9?�8h�\?n?�?�?�?��? _S����  �Aa{p���m�Y_�Ed�� T=�nD4vnCIO�䑎II@`�O��_�OP�E�C.r��WP�OWE	�� �X@�f��$�$Cd�S����i��A3�3� �@��SI��G�P0�QIRT�UAL�O
QAAV�M_WRK 2 �7U 0  �5Q�n_zXk_�] ��\	�P�]�_3�8P��_�_�Ve�\#m/o��Q5ojo|o�dHPBS��� 1Y� <Xo�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯�ݯ�bC$�AXLM��@���c  �d�IN����P+RE
�E�J�-�'_UP��[�7QHP?IOCNV_��k �	�Pr�US>��g�cIO)�V 1]U[P $E`��Q0ս9lҿ8P?�� � ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o�o�o�o�m�LAR�MRECOV �a��-���LMD/G ��ɰ��LM_IF  ���ை����z�v���%�6�, 
 6�_��r� ��������̍$w��� ׏��8�J�\�n�����NGTOL  �a� 	 A �  ��ț�PPI�NFO ={� <v����1��  I�3�a�"rP��� t��������ί���>�o����j�|��� ����Ŀֿ������0�B�PzPPLIC�ATION ?����+��HandlingTool ��� 
V9.30�P/04ǐM�
�88340�å�F90����202�ť�|�Ϭ�7DF3���M̎�NoneM��FRAM� �6��Z�_ACTI�VE�b  sï� � p�UTOMO�Dz�A���m�CH�GAPONL�� ���OUPLEDw 1ey� �������g�CURE�Q 1	e{  T*���	p��xw���#r�g���e�HN����{�HTTHK)Y��$r��\[�m� ���O�	�'�-�?�Q� c�u����������� ��#);M_q ������ %7I[m� ��/���/!/ 3/E/W/i/{/�/�/�/ ?�/�/�/??/?A? S?e?w?�?�?�?O�? �?�?OO+O=OOOaO sO�O�O�O_�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q��c���1�TO��|��p�DO_CLEA�N��n��NM  �� �B�T��f�x���%�DSPDgRYR��m�HI���@/�����,�>� P�b�t���������ίj�MAXa�ۄ�������Xۄ������p�PLUGG��܇�Ӯ��PRC��B�" ��ׯF�OK���^ȔSEGF��K�� �����.�����,�8>�v���LAPӟ� ��Ϥ϶��������π�"�4�F�X�j߯�T�OTAL�7���U�SENUӰ�� ����ߖ�1�RGDI_SPMMC����C����@@Ȓ��O�ѐ�����_STRING 1
�ۿ
�M��S�l�
A�_ITE;M1K�  nl�g� y������������ 	��-�?�Q�c�u����������I/O SIGNALE��Tryout� ModeL�I�np��Simul�atedP�Ou�tOVER�RА = 100�O�In cyc�lP�Prog� AborP�~��StatusN��	Heartbe�atJ�MH F�aul��Aler�	�������*<N`  ׃G�ׁY�c��� ��////A/S/e/ w/�/�/�/�/�/�/�/wWOR��G�-1� ?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO�cOuO�O�O�NPO E��@E;�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8oJo�BDEV�Nu`�O bo�o�o�o�o�o�o ,>Pbt�������PALT��E?�A�S� e�w���������я� ����+�=�O�a�s����GRI�G뽑 1������	��-�?� Q�c�u���������ϯ�����)�����R �a�՟;��������� ѿ�����+�=�O� a�sυϗϩϻ���O�PREG��y��� -�?�Q�c�u߇ߙ߫� ����������)�;��M�_�q����$AR�G_-0D ?	��������  	$���	[��]���������SBN_CONFIG���� ��CII�_SAVE  ���)���TCEL�LSETUP ���%  OME�_IO����%M�OV_Hn�����R�EPd�����UTO/BACKY���#�FRA:\��� ����)�'`rl ��&� 7�"� 24�/06{  09:_35:24������͓����� �+=Oas��������� �/1/C/U/g/y/�/ /�/�/�/�/�/	?�/ -???Q?c?u?�?�?p�ׁ  _��_\�ATBCKCTL.TM���?�?�?O\ O��INI�Y��-���MESSA�G9�GA)��RKODGE_Ds�<��zH�Ow`�O��PAUS��@ !��� ,,		�����O �G�O__#_%_7_q_ [_�__�_�_�_�_�_��_%o���D�@TSK  �M&,O���UPDT�@EGd��`�FXWZD_E�NBED��fSTApDE��e��XIS�?UNT 2��&��(�� 	\` ��� �� ���$ N`� ���  i�b	��\b�p�p�<��� �Ug~pj3N� �rZ�l�o��W�IPb�D$��yk~����dMETc�2�LfE� P qA�pA�G�AD��sB S8A��BR�o�}>�Ì�?R=a?���@5��?7g�@`��}�SCRDCFG �1�� 	�A�&������ ԏ�����Q=��� H�Z�l�~�����	�Ɵ -����� �2�D���域���GR�`�`�O����0NA����	���_EDC@1�n�� 
 �%{-�0EDT-q�0���%�p��"���Q-���������x����  ����!2����*�RIE����*�q���ϧ���3 bϮ�@Ͻϯd?����� =�O���sϏ�4.ߞ� {�����W���	�߱�?ߏ�5��j�G���΀#������}�6 ��6��Z�����Z�����I��7����� &��λ�&m����B��8^ҿ�����̀��9K�o��9*�w����S�`�;��CR�� ��B/T//�/���w//��РNO_D�EL����GE_U�NUSE���IG�ALLOW 1���   (�*SYSTEM*��s	$SERV�_GR�;B0�@RE�GK5$m3�|B0N�UMp:�3�=PM�U� �uLAY��p�|PMP�ALD@�5CYC1�0�.�>�0�>CULSU�?�=�2�AM3�LOWDBOXO{RIt5CUR_D@~�=PMCNV�6�D@10�>�@T�4DLI�`=O_9	*PROGRAJ4PG_MI�>��OPAL�E_U�PB7_B>$FLUI_RESU�70p_z?�_�TMRY>h0�,�/�b�_�_o o 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����������"LAL_?OUT 1;l����WD_ABOR��0?d�ITR_R_TN  ����~g�NONSTOǠ��� 8CE_R�IA_I0���ۀ��ŀFCFG� ��۔��_�LIMY22ګ� �  � 	�i�J��<e�g��5��P� 9�������
���u��PA�QPGP 1�����Q�c�u�4��CK0����C1��9ҭ�@���PC��CV���]��d��l��s����0���C[٤m���v���������� C����-����?�ÂHE� O�NFI�Pq�G�G_�P�@1�  �%�������ǿٿ�����G�KPAUSfaA1�ۃ �2 �W��Eσ�iϓϹ� �����������#�I�@/�m��eߣ��M���NFO 1"��� �7��ߖ���³��A����/^$C3������BL�� =�<��Į�4l���A�؏C�3�E�ŀO��c�CO�LLECT_�0"�[�����EN�@���y���k�NDE���"�3�"12�34567890���\1�� ��֕H&��)M�r�\,L�^� ��]+������������ C 2�Vhz ������
 c.@R�v���������� �����IO !���q���u/�/�/l�/C'TR�2"'-�(�P^)
��.R��#R-�*W� 9_MO5R�$� �;�l5 ��l9�?r?�?�?�?�;�E2��%S=,W�?$@�@��C�PK)DցC�R�&u�XOWA~WBC4  A�q����Px�PA"@C�z  B�@CG�B|8��AC  @yB���Pց:d��43 <#�
@�E���I�O�C=AI��%'GM?�C�(S=����Qd=AT_DEF�PROG �;%��/m_APINUS�E�V�ۅ�TKEY?_TBL  s�ہ����	
��� !"#$%&�'()*+,-.�/�:;<=>?�@ABCDPGHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������Ga��͓���������������������������������耇�������������������s��!�PLCK�\8���P�PSTAn��T�_AUTO_DOr��NFsIND��<�n��R_T1w�T2N����5ŀT{RLCPLETE����z_SCREE�N �k�cscÂU��MM�ENU 1)O� <�[_#�q��,� a���>�d���t���ӏ ����	�����Q�(� :���^�p�������̟ �ܟ�;��$�q�H� Z����������Ưد %����4�m�D�V��� z���ٿ��¿�!��� 
�W�.�@ύ�d�vϜ� �ϬϾ������A�� *�P߉�`�r߿ߖߨ� �������=��&�s� J�\������������'�,�p_MANgUAL�EqDB
1�2�v�iDBG_E7RRLIP*�{h!� 0�������~g�NUMLIM�s�:QOE�@DBPXWORK 1+�{��>Pbt��-�DBTB_�q Q,��kC3!VD!DB_AWAYo�h!GCP OB=9��A�_AL���o��k�Y�p�uO@`�_��� 1-�+@
�-k-6[��_M&+pIS�`�@"@��ONTIM�w�&OD��&
�U;MOTNEND�_�:RECORD ;13�{ ��[CG�O�f!T/[K� �/�/�/�/_(�/�/f/ ?�/??Q?c?�/?�? ?�?,?�?�?OO�? ;O�?_O�?�O�O�O�O (O�OLO_pO%_7_I_ [_�O_�O�__�_�_ �_�_l_!o�_,o�_io {o�o�oo�o2o�oVo /A�oeP^ �
���R�� �=��a�s������ ��*�ߏN���'��� ԏ]�̏��������ɟ ۟v���n�#���G�Y��k�}���TOLEoRENC�B�0�� L��g�CSS�_CNSTCY +24	�t���.������0�>�P� b�x���������ο�����(�:�äDEVICE 25ӫ ��ϟϱ��� ��������/�Aߟ�ģHNDGD 6ӫ� CzT�.!ơ_LS 27t�S� ����������/�U��ŢPARAM �8Gb�A�Ք�R�BT 2:�8�<���Ck�A� ·�  � A���.�SB���A�B�O  ���������.�� �,���A�A�C�����c�u����C�A�D���k�pz�A,�A��HA�c��A� 	�?(uL^p����A�Bt/��D��C��_ �	 A=��A�BffA#33A}Ҋ���A�A�Cf��a��A��J��7B]��B���BffB}ᴠ�33C$.@R� ( �� �A����
/�� //)/;/�/_/q/�/ �/�/�/�/�/�/<?? %?r?I?[?m??�?�? �?�?�?&O8O�PObO MO�OqO�O�O�O�O�O _�OOL_#_5_�_ Y_k_�_�_�_�_ o�_ �_6oooloCoUogo �o�o�o�o�o�o �o 	h�O�w�� ���
��.�	__ I'�1_�q������� �ˏݏ���%�r� I�[����������ǟ ٟ&����\�3�E�W� ���ȯ���ׯ�"� �F�1�j�E�s����� m�������ѿ�0�� �f�=�O�a�sυϗ� �ϻ��������'� 9�Kߘ�o߁�����[� ���(��L�7�p�� m����������� $�����l�C�U��� y����������� �� 	V-?�cu� ���
��@+ dO�s���� ����*///`/7/ I/[/m//�/�/�/�/ ?�/�/?!?3?E?�? i?{?�?�?�?�?�?�? �?FO�jOUOgO�O�O �O�O�O�O__�'O 9OO=_O_�_s_�_�_ �_�_�_�_�_oPo'o 9o�o]ooo�o�o�o�o �o�o:#5� �O����� ���$��H�Fz�$DC�SS_SLAVE ;���w���`�_4�D  w���AR�_MENU <w� >�؏���� �2�^rǏ\�n�\���SHOW 2=w� � fr[q�� ��Ə�����,�>�D�b�t��� ����ҟ ϯ����)�P�M� _�q���������˿ݿ ���:�7�I�[ς� |Ϧ��ϵ��������� $�!�3�E�l�fߐύ� �߱���������� /�V�P�z�w���� ����������@�:� d�a�s����������� \���*�H�N�K] o�������� 28�GYk} ������" �1/C/U/g/y/�/� �/�/�/��//?-? ??Q?c?u?�/�?�?�? �/�??OO)O;OMO _O�?�O�O�O�?�O�? �O__%_7_I_pOm_ _�_�O�_�O�_�_�_ o!o3oZ_Woio{o�_ �o�_�o�o�o�o Do-Se�o��o� �����.�=��O���CFG >Ɨ����q��d�MC:\��L%04d.CSV\�Ҁpc�������A ՃCH݀z�v�w(�#��q���:��J�8�7���JP�(j�)�́�p+�n��RC_OUT -?z�����a��_C_FSI ?���  |�����@�;�M� _���������Я˯ݯ ���%�7�`�[�m� �������ǿ���� �8�3�E�Wπ�{ύ� ������������� /�X�S�e�wߠߛ߭� ���������0�+�=� O�x�s�������� �����'�P�K�]� o��������������� ��(#5Gpk} ����� � HCUg��� ����� //-/ ?/h/c/u/�/�/�/�/ �/�/�/??@?;?M? _?�?�?�?�?�?�?�? �?OO%O7O`O[OmO O�O�O�O�O�O�O�O _8_3_E_W_�_{_�_ �_�_�_�_�_ooo /oXoSoeowo�o�o�o �o�o�o�o0+= Oxs����� ����'�P�K�]� o�����������ۏ� ��(�#�5�G�p�k�}� ������şן ���� �H�C�U�g������� ��دӯ��� ��-� ?�h�c�u��������� Ͽ�����@�;�M� _ψσϕϧ������� ����%�7�`�[�m� ߨߣߵ��������� �8�3�E�W��{�� ������������� /�X�S�e�w������� ��������0+= Oxs����� �'PK] o������� �(/#/5/G/p/k/}/ �/�/�/�/�/ ?�/?�?H?C?U3�$DC�S_C_FSO �?����1� P  [?U?�?�?�?�?�?O 
OO.OWOROdOvO�O �O�O�O�O�O�O_/_ *_<_N_w_r_�_�_�_ �_�_�_ooo&oOo Jo\ono�o�o�o�o�o �o�o�o'"4Fo j|������ ���G�B�T�f��� ������׏ҏ���� �,�>�g�b�t����� ����Ο�����?� :�L�^���������ϯ�ʯܯg?C_RPI~>�?�;�d�_�
��}?.�p����ݿj>SL�@���9�b�]� oρϪϥϷ������� ���:�5�G�Y߂�}� �ߡ����������� �1�Z�U�g�y��� ����������	�2�-� ?�Q�z�u��������� ����
)RM _q������ �*%7Irm �����/� ϛ�,�/W/�/{/�/ �/�/�/�/�/??? /?X?S?e?w?�?�?�? �?�?�?�?O0O+O=O OOxOsO�O�O�O�O�O �O___'_P_K_]_ o_�_�_�_�_�_�_�_ �_(o#o5oGopoko}o �o�o�o�o�o �o HCUg��� ����� �����NOCODE }@������PRE_CHK �B��3�A 3��< �7�🵧����� 	 < �����?#ۏ%�7�� [�m�G�Y�������ٟ �ş�!����W�i� C�����y�ïկˏ�� ����A�S�-�_��� c�u���ѿ������ �=��)�sυ�_ϩ� �ϕ��������'�9� ��E�o�I�[ߥ߷ߑ� ��������#����Y� k�E���{����� ������C�U��=� ����w���������	 ����?Q+u�a ������) ;_qg�Y�� S����%/�/ [/m/G/�/�/}/�/�/ �/�/?!?�/E?W?1? c?�?���?�?o?�? O�?�?AOSO-OwO�O cO�O�O�O�O�O_�O +_=__I_s_M___�_ �_�_�_�_�?�_'o9o o]oooIo�o�oo�o �o�o�o#�oGY 3E��{��� ��o�C�U��y� ��e�����������	� �-�?��K�u�O�a� ��������͟��)� �1�_�q��}����� ��ݯ�ɯ�%���1� [�5�G�����}�ǿٿ �������E�W�1� {ύ�G�u����ϯ��� ���/�A��-�w߉� c߭߿ߙ��������� +�=��a�s�M��� �ϑ�������'�� 3�]�7�I�������� ����������GY 3}�i������ ��C/y �e������ �-/?//c/u/O/�/ �/�/�/�/�/�/?)? �?_?q?K?�?�?�? �?�?�?�?O%O�?IO [O5OO�OkO}O�O�O �O�O_�O3_E_;?-_ {_�_'_�_�_�_�_�_ �_�_/oAooeowoQo �o�o�o�o�o�o�o +7aW_i_�� C�����'�� K�]�7�i���m��ɏ ۏ�������G�!� 3�}���i���ş�� ����1�C��g�y� S�e����������ѯ �-���c�u�O��� ����Ͽ�ןɿ�)� ÿM�_�9�kϕ�oρ� ���Ϸ������I� #�5�ߑ�kߵ��ߡ� ������3�E���Q� {�U�g��������� ���/�	��e�w�Q� �������������� +Oa�I�� ����� K]7��m�� ���/�5/G/!/ k/}/se/�/�/_/�/ �/�/?1???g?y? S?�?�?�?�?�?�?�? O-OOQOcO=OoO�O �/�/�O�O{O�O_�O _M___9_�_�_o_�_ �_�_�_oo�_7oIo #oUooYoko�o�o�o �o�o�O�o3Ei {U������ ��/�	�S�e�?�Q� ������я㏽��� �O�a�������q� ��͟�������9� K�%�W���[�m���ɯ �����ٯ�5�+�=� k�}����������� ��տ�1��=�g�A� Sϝϯω����Ͽ��������Q�c�����$DCS_SGN� CS����#�M�14-�JUN-24 0�9:43 E��06��39������� X�L�������������Д���M��Þ�ǧj�����{�VE�RSION ���V4.2.�10�EFLOG�IC 1DS���  	�D���X�k�X�z�M�P�ROG_ENB � ��b��Л�U?LSE  ����M�_ACCLI�M��������WRSTJNT�����w�EMO���ѷ�L��INIOT EZ�O���OPT_SL ?�	S�1�
 	�R575�Ӆ�74*��6��7��5A��1��2��l���G�h�TO  t���.�H�V?�DEX��d����FPATHw A��A\4����HCP_CLNTID ?+�b� l������IAG_GRP� 2JS�� �a[��D�  D�� �D  B�  ;B�@ff��/CB�@[��W�@��q��B�N��C�-Bz�w�Bp@e`���mp3m7 �78901234�56�*�[�� � Ao�mAj�1AdA]��
AW|�AP��AJ-AC�/A;�A4�H���@�  Aʩ�A�A3!_A�@@��B4��� ��t���
�u�ƨApffAj��yAeK�A_��AY��AS�� MC�AF��A@ �O�+/=/O$�O�c K�w(@�X�?8��@��y�/�/�/�/�/8��;d�2�5?@~�ff@x1'@q���@kC�@d��D@]��@Vv�6?H?Z?l?~?8�s�0l��@e���@^��@W\)@O��@H�0�?<@7K�@.V��?�?�?�?
O8S�@M00G<@A���@<1@5���@/l�@(�Ĝ@!�0�\ NO`OrO�O�Ox'g�L_ K�;_�_�__g_�_�_ �_�_o�_�_�_Yoko@Io�o�o+o�oX�"�� 2�17A�@J>���R
q?�33?wY��r��J�7'Ŭ2q63p4w�F>r��LJ�@�p�Zr�
=�@�@�Q�jq��@G Ah�@���@�T= c<���]>*�H>�V>�3�>����J<���C<�p�q�x��� ��?� �C� � <(�U�� 4Vr�33��@
���A@��?R�oD� �mR�x���Q��t�����Z�Џ��؏�,��i?��7N�>�(�y>�@Z�=���Jo��G�v�G�J �B�E�����a��@ǐ�@���@��@OQ�?L ���ŲI�P���&�
��'��@�K�����Ag�q�PC�  ?C���Cuy�
����ʯ ?տNL��>�;����B�?� >穪��*���
��S������F�ĺ��/��H��>(���P4���X��v����*
���A�?�EC�gF�ǿ B��ֿ����E�Tt���X�!�AB�І��fzWC� 
éF�
��Iϗ�CT_CONFIG Ky3���e���B�STBF_TTS��
����"���t����{�MAU�����MSW_CF���L  K �O�CVIEW	�MI�U����߭߿� ���������0�B� T�f�x�������� ������,�>�P�b� t�������������� ��(:L^p� �����  �6HZl~�������/��R%CB�N��!�X. F/{/j/�/�/�/�/�/���SBL_FAULT O9*^�1GPMSK��7���TDIAG PԺ�U����q�UD1: 67�89012345 q2�q���%P�ϭ? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �a6�I'�
�?_�ƟTRECPJ?\:
 j4\_�7u[�?�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�O�O�_ _�UMP_OPTION��>q�TRB���9;uP�ME��.Y_TE�MP  È�g3B����p�A�pytUNI'��ŏq6��YN_BRK �Qt�_�EDITO�R q&qh�r_2PE�NT 1R9) � ,&MAI�N A_BARR�A�P�p  ?&SEGU*�'���.&COLOC�A_PRENSA� VIS$r��t��x�BASE_IR�����&PIC�K1_PLACE�0Z��&ЁU�P~�ޏ�&
P�EGA_�pNO ��.���p���U�-��;���&(�S�E?STEIRAf�L��ւR������&SUMIRZ���p����a�����[��0���p�#��/�������ï���ί�� ��A�(�e�w�Jq�p�MGDI_STA�u~��q�uNC_I?NFO 1SI��b�������Կ�쮳��1TI� �P�o#��G�
G�d�o }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߯���������Hu�  �2�D�R�j�R�x�� ������������� ,�>�P�b�t������� ������Z��#5 Ga�k}���� ���1CU gy������ ��	//-/?/Yc/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?��?O%O 7OQ/GOmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �?Ooo/o�_[Oeo wo�o�o�o�o�o�o�o +=Oas� �����_�_�� '�9�So]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�K�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�C�5�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ��������!�;�M� W�i�{�������� ������/�A�S�e� w��������������� +E�Oas� ������ '9K]o��� �1����/#/= G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?��? �?	OO5/?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�?�_�_oo-O #oIo[omoo�o�o�o �o�o�o�o!3E Wi{����_�_ ����7oA�S�e� w���������я��� ��+�=�O�a�s��� ������ߟ��� /�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������͟ ׿����'�1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߫�ſ������� ��;�M�_�q��� �����������%� 7�I�[�m�������� ���������)�3E Wi{����� ��/ASe w��������� /!+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?/ ��?�?�?�?/#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�?�_�_�_ �_Oo-o?oQocouo �o�o�o�o�o�o�o );M_q�� �_����	o�%� 7�I�[�m�������� Ǐُ����!�3�E� W�i�{�����ß՟ 矝���/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߩ����� �������1�C�U� g�y���������� ��	��-�?�Q�c�u� ���߫����������� );M_q�� �����% 7I[m���� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?���?�?�?�?� OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�?�?�_ �_�_�_�?�_o#o5o GoYoko}o�o�o�o�o �o�o�o1CU gy�_�����_ �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q��y� ����˟�۟��%� 7�I�[�m�������� ǯٯ����!�3�E��W�i��� �$EN�ETMODE 1�U�� W ���������»��RROR_PROG %���%�����TAB_LE  ����Q�c�uσ��SEV�_NUM ��  �������_AUTO_EN�B  ̵��ݴ_;NO�� V����}��  *���������������+����(�:���FLT9R����HIS�Ð������_ALM 1]W�� �������+;����������0�?�_����  �����²u꒰T�CP_VER �!��!��@�$EX�TLOG_REQ�v������SIZ\����STK��������TOL  ���Dz~��A= ��_BWDU�*�Z�V�ǲ?�DID� ;X�Z���<��[�STEPl�~�|����OP_DO����FACTORY�_TUNv�d��D�R_GRP 1Y��`�d 	p�.°� �*u����RHB ���2 ��� �e9 ���bt�� B��!C'��CۺDC���#C��D!�v�A���B�&�B=�A���A���BLZ������
C.gR  A�A">A.�@"�?�Βu
 I�������<��n���_/�(/�	�  �F!A�  @�3�3R"�33�@UUTn*@P  /ȷ�>u.�>*���<��ǊE��� F@ �"�5�W�%�J��NJ�k�I'PKH�u��IP�sF�!���?�  �?�/9�<9��896C�'6<,5����.� R�D��"� ��t� 	q4 "�ơ���EATUROE Z�V�Ʊ�Handl�ingTool ��5��Engl�ish Dict�ionary�74�D St�0ard��6�5Analog� I/O�7�7gle Shift O�uto Soft�ware Upd�ate%Imati�c Backup��9SAground� Edit�0�7C_amera�0F�?�CnrRndIm�XC�Lommon �calib UI�C�FnqA�@Monoitor�Ktr�0?Reliab@�8�DHCP�IZat�a Acquis��CYiagnos�OA�1[ocume�nt Viewe��BWual Ch�eck Safe�ty�A�6hanc�ed�F�:�UsnPF�r�@�7xt. D7IO �@fiRT�Wwend�PErr�@QLQR�]�Ws�Yr�0��P E�:FCTN_ Menu�Pv S�8gTP In'`f�acNe�5GigE�`nrej@p Mas_k Exc�Pg�W�HT^`Proxy� SvoT�figh�-Spe�PSki�D�eJP�Pmmun�icN@ons�hu�rE`'`_�1abconnect 2x�ncr``struH�2z>peeQPJQU��4KAREL C�md. L�`ua��husRun-Ti��PEnvkx(`el� +R@sP@S/W��7License��Sn\�PBook(System)�:MACROs,�b?/Offse@�uaH�P8@_�pMR�@��BP^MechSt�op�at.p6R�ui�RKj�x�P�0P@)��od@witchȘ�>�EQ.���Op�tmЏ>��`fil�n\=�gw�uult�i-T�`tC�9PC�M funHwF�o�3T�R?�f�Regi��pr�`I�rigPF�V����0Num S�elb����P Ad�ju�`���J�t�atu��
�iZ�5R�DM Robot>�0scove�1F��ea7��PFreq� Anly�gRe�m`��Qn�7F�R�S�ervo�P���8S�NPX b�rNSN^`ClifQɮB�Libr�3鯢0 �q�����o�ptE`sGsag?��4�� -C���;��/I_mB�M�ILIBk�E�P OFirm6BU�PEc�Acck@sKTPT9X_C�eln����F��1�V�orqu>@imula�A�A�u��Pa�qU�j@t�Ã&�`ev.B��.@riP޿USB port �@�iP�PagP��R �EVNT�ϗ�nexcept�P��t�X�ſX�]VC�Ar�b�bf�V2PҦ�$�����SܠSCصV�S�GEk�a�UI�;Web Pl!��ާ���Խ`�TeQfZD?T Appl�d�:x�ƺ� �GridV�play�R�WD4�R
�.�:n�EQ+��r�-10iA/7L�*��1Graphi�c���5dv�SDC�SJ�ck�q�5la�rm Cause�/��ed�8Asc�ii�a��Load�nP�Upl,�Ol�0�AGu�6N�`���yFyc@�r�����P�V��Jo��m� c��R���c���m�./������Q�2*u:eRA`J��P�ٶ4eqinL�����8NRT��9O}n�0e Hel�H�J�`oI�allet�iz?�H�����_�t�r�[ROS Eth�q��T@e�ׅ�!��n�%�2D�tPkgp&Upg~��(2DV-�3D� Tri-jQEA�ưDef.qEBa)pdei��� �b�ImπF�f��n�sp.q=�464M?B DRAMZ,#�FRO5/@ell��<�Mshf!r/�'c�%3@pLƖ,ty�@s˒xG��m��. [�� ��BU���Q�B�=mai�P߫�]hQ����@q6wlu��H��^`�xR�?eL� Sup������0�P�`cr��@�R���b�x���pr1uest�Crt~QQ��ߋL!��4O��q$�K��l� Bui7�n��A'PLCOO�EVl%��sCGU�OCRG�Ob��DR��O
TLS_&��BU/_��K�qN_&d�TA�OxVB�_�Wp�ܑZ���_TCB�_ �V�_�W���WF+o�V��O�W._�W�ņoTE�H�o�f�O�gt�oT	Ej�xVF�_w�_xV�GoTwBTw~oxVH�xVIA��v�xVLN�yUMz�boH�f_xVN�xVP�H��^xVR&xVS��܇ʏ��W��v���gVGF:�L�P2_�h��h�V�h��_g�D���h�FFoh��g�R�D�� TUT��0�1:�L�2V�L�TB�GG��v�rain�UI��
%HMI���pon��m��f�"�F�&K�AREL9� �TP�j��<6 SWIM7ESTڢF0O�<5�
"a�X�j������� ͿĿֿ���'��0� ]�T�fϓϊϜ����� ������#��,�Y�P� bߏ߆ߘ��߼����� ����(�U�L�^�� ������������� �$�Q�H�Z���~��� ����������  MDV�z��� ���
I@ Rv����� �///E/</N/{/ r/�/�/�/�/�/�/? ??A?8?J?w?n?�? �?�?�?�?�?O�?O =O4OFOsOjO|O�O�O �O�O�O_�O_9_0_ B_o_f_x_�_�_�_�_ �_�_�_o5o,o>oko boto�o�o�o�o�o�o �o1(:g^p ������� � -�$�6�c�Z�l����� ����Ə����)� � 2�_�V�h��������� ����%��.�[� R�d������������ ���!��*�W�N�`� �����������޿� ��&�S�J�\ωπ� �Ϥ϶��������� "�O�F�X߅�|ߎߠ� �����������K� B�T��x������ �������G�>�P� }�t������������� C:Lyp ������	  ?6Hul~� ����/�/;/ 2/D/q/h/z/�/�/�/ �/�/?�/
?7?.?@? m?d?v?�?�?�?�?�? �?�?O3O*O<OiO`O rO�O�O�O�O�O�O�O _/_&_8_e_\_n_�_ �_�_�_�_�_�_�_+o "o4oaoXojo|o�o�o �o�o�o�o�o'0 ]Tfx���� ���#��,�Y�P� b�t������������ ���(�U�L�^�p� ���������ܟ�� �$�Q�H�Z�l�~��� �����د��� ��M�D�V�h���  H552}�v��21��R78��{50��J614���ATUPͶ545z͸6��VCAM��wCRI�UIFͷ�28	�NRE��5�2��R63��SC�H��DOCV]�C�SU��869ͷ0^ضEIOC9�4���R69��ESET����J7��R68޴�MASK��PR�XY!�7��OCOB��3帨���̸3�[J6˸53��H2��LCH��OPLGz�0�MHCR��]S{�MCS�0��{55ضMDSW��v�OP�MPR�tM�@�0̶PCM ƃR0���ض��@�5�1�51<�0�P�RS��69�FR�D�FREQ��M�CN��93̶SN�BAE�3�SHLB���M��M���2̶H{TC�TMIL����TPA��TPT�X��EL��Ѐ�8�������J95,�T�UT�95�UE�V��UEC��UF]R�VCC��O��wVIP�CSC,��CSG8�r�I��W�EB�HTT�R�6C�N�CGIG���IPGS)RCv�DG�H77���6ضR85��R6�6�R7��R:�R[530�680�2�Rq�J��H�6<�6,�QRJح�0�4�6o�64\�5�NVDv��R6��R84Thg����8�90\�6��J93�91� �7+���,�D0oF��CLI���CMqS�� �STY���TO�q���7�N]N�ORS��J% ���j�OL(END굶L��Sf(FVRΘ�V3D���PB�V,�APL��AP�V�CCG�CC�R|�CD��CDL�@CSBt�CSKv��CT�CTBL9���U0,(C��y0L8C���TC �y0�'TCv(7TC��CTE\ƌ�07TEh��0��TUFd8F,(GL8GI
�8H�8I��E@�87�WCTM,(M�8M@8UN�8PHHPL8Rd8�(TSd8W�I@V�GF�GP2��P2p���@�H{7VPD�H�F �VPSGVPRƘ&VT��YP��VT�B7Vs�IH��VXI aH'VK��VGene�����_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A� S�e�w���������џ �����+�=�O�a� s���������ͯ߯� ��'�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a?�s?�?  H55hT�1�1[U�3�R78�<50�9Jw614�9ATU�T��4545�<6�9VsCA�D�3CRI,K�UI8T�528-JN�RE�:52JR6�3�;SCH�9DO�CV�JCU�486u9�;0�:EIO�T�sE4�:R69JEgSET�;KJ7K�R68�JMASK^�9PRXYML7�:OCO\3�<�J)P��<3|ZJ6�<53��JH�\LCH\ZO�PLG�;0�ZMH�CR]ZSkMCS��<0,[55�:MD�SW}k�[OP�[M�PR�Z�@�\0�:PCMLJR0�k)P�:l)`�[51K51|�0JPRS[69�|ZFRD<JFRE�Q�:MCN�:93��:SNBA}K�[SHLB�zM�{�@ll�2�:HTC�:TMsIL�<�JTPA�JoTPTX�EL�z�)`�K8�;�0�JJ9�5\JTUT�[95�|ZUEVZUEC�\ZUFR<JVCC���O<jVIP,�C;SC\�CSGlJ�@�I�9WEB�:HT�T�:R6{L��CG�{�IG[�IPGS���RC,�DG�[H�77�<6�:R85n�JR66JR7[�R|R53{68�|2�Z�@Jml,|6�|6\JR�\	P|4ZL�6�64��5�k�NVDZR6+kRC84<���IP,�8���90���KJ9�\9�1��̫7[KIP\JDu0�F��CLI�l�KCMS�J9��:STY,�TO�:�@�K�7�LNN|ZORSb<jJ��MZZ|OLK�WEND�:L�S��wFVR�JV3D,��KKPBV\�APL��JAPV�ZCCGn�:CCRjCD�wCDL̚CSB�J�CSK�jCTK�CCTB��\���\�C�z4���CL�TCLJ�l�TC��TCZCcTE�J��|�TE�J���<�TF��F\�GR��G��l�Hl�I�z�)�l�k�CTM\�M�\�M��Nl�P,�P���R��;�TS��W���̚VGF��P2���P2�z �VkPDFLJVP;�7VPR��VT�;� ��JVTB��V�KI�H�VِM�<�VKz,�V{�Gene�8 �83EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w��������� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y������� ��������	-? Qcu����� ��);M_ q������� //%/7/I/[/m// �/�/�/�/�/�/�/?�!?3?E?W?i?{?�7��0STD�4LANG�4�9�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D��V�RBT�6OPTNm��������Ǐُ ����!�3�E�W�i��{�������ß�5DPN�4�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߡ���ted �4�8�� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯٯ������*�<�pN�`�r���99����$FEAT_A�DD ?	��������  	��ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?Q�cu�����DE�MO Z��   ���}�� '��0�]�T�f����� ����������#�� ,�Y�P�b��������� ��������(�U� L�^������������ ܯ���$�Q�H�Z� ��~��������ؿ� �� �M�D�Vσ�z� �Ϧϰ��������
� �I�@�R��v߈ߢ� �����������E� <�N�{�r������ �������A�8�J� w�n������������� ��=4Fsj |������ 90Bofx� ������/5/ ,/>/k/b/t/�/�/�/ �/�/�/�/?1?(?:? g?^?p?�?�?�?�?�? �?�? O-O$O6OcOZO lO�O�O�O�O�O�O�O �O)_ _2___V_h_�_ �_�_�_�_�_�_�_%o o.o[oRodo~o�o�o �o�o�o�o�o!* WN`z���� �����&�S�J� \�v����������ڏ ���"�O�F�X�r� |�������ߟ֟�� ��K�B�T�n�x��� ����ۯү���� G�>�P�j�t������� ׿ο����C�:� L�f�pϝϔϦ����� ��	� ��?�6�H�b� lߙߐߢ�������� ���;�2�D�^�h�� ������������
� 7�.�@�Z�d������� ����������3* <V`����� ���/&8R \������� ��+/"/4/N/X/�/ |/�/�/�/�/�/�/�/ '??0?J?T?�?x?�? �?�?�?�?�?�?#OO ,OFOPO}OtO�O�O�O �O�O�O�O__(_B_ L_y_p_�_�_�_�_�_ �_�_oo$o>oHouo lo~o�o�o�o�o�o�o  :Dqhz �������
� �6�@�m�d�v����� ��ُЏ����2� <�i�`�r�������՟ ̟ޟ���.�8�e� \�n�������ѯȯگ ����*�4�a�X�j� ������ͿĿֿ��� �&�0�]�T�fϓϊ� �������������"� ,�Y�P�bߏ߆ߘ��� ����������(�U� L�^��������� ���� ��$�Q�H�Z� ��~������������� �� MDV�z ������� I@Rv�� �����//E/ </N/{/r/�/�/�/�/ �/�/�/
??A?8?J? w?n?�?�?�?�?�?�? �?OO=O4OFOsOjO |O�O�O�O�O�O�O_ _9_0_B_o_f_x_�_ �_�_�_�_�_�_o5o ,o>okoboto�o�o�o �o�o�o�o1(: g^p����� �� �-�$�6�c�Z� l�������ϏƏ؏� ��)� �2�_�V�h��� ����˟ԟ���%� �.�[�R�d������� ǯ��Я���!��*� W�N�`�������ÿ�� ̿����&�S�J� \ωπϒϿ϶����� ����"�O�F�X߅� |ߎ߻߲�������� ��K�B�T��x�� ������������ G�>�P�}�t�������>��  ���� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t��������� ο����(�:�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz�����y  �x�q���&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p������q�p�x�� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p���������������$FEA�T_DEMOIN�  �� ������INDEX����ILE�COMP [w���B���8 SETUP2� \BL��  N w5_�AP2BCK 1�]B	  �)�����%���� E �	���5�Y �f��B�� x/�1/C/�g/� �/�/,/�/P/�/t/�/ ?�/??�/c?u??�? (?�?�?^?�?�?O)O �?MO�?qO O~O�O6O �OZO�O_�O%_�OI_ [_�O__�_�_D_�_ h_�_�_
o3o�_Wo�_ {o�oo�o@o�o�ovo �o/A�oe�o� ��N�r�� �=��a�s����&� ��͏\�񏀏���"� K�ڏo�������4�ɟ X������#���G�Y� �}����0���ׯQ	�� P� 2� �*.VRޯ(���*+�Q���W�{�e���PC������FR6:��ؾg�����T   �2����\� x��d�*.F�D�ϕ�	ó����o�ߓ�STM�9����ư%�d��ψߓ�H U߻�Jש�f�x���GIF�A�L�-���8�ߑ��JPG�����Lձ�n�����JS��H�����6���%�
JavaScrgiptt���CSe����Kֹ�v� %C�ascading� Style S�heets��j�
�ARGNAME.SDT'��O�\;���[�k|(k DISP*rUOп���� �
TP�EINS.XML�/�:\CcC�ustom To�olbar��	PASSWORD�~��FRS:\��� %Pass�word Config/c�Q/�J/ �/���/:/�/�/p/? �/)?;?�/_?�/�?? $?�?H?�?l?�?O�? 7O�?[OmO�?�O O�O �OVO�OzO_�O�OE_ �Oi_�Ob_�_._�_R_ �_�_�_o�_AoSo�_ woo�o*o<o�o`o�o �o�o+�oO�os� �8��n�� '���]�����z� ��F�ۏj������5� ďY�k��������B� T��x�����C�ҟ g�������,���P�� �������?�ί�u� ���(���Ͽ^�󿂿 �)ϸ�M�ܿqσ�� ��6���Z�l�ߐ�%� ���[����ߣߵ� D���h�����3��� W����ߍ���@�� ��v����/�A���e� �����*���N���r� ����=��6s �&��\�� '�K�o�� 4�X���#/� G/Y/�}//�/�/B/ �/f/�/�/�/1?�/U? �/N?�??�?>?�?�? t?	O�?-O?O�?cO�?��OO(O�O�F�$F�ILE_DGBCK 1]���@��� �< �)
SUMMARY.DG�O�sLMD:�O;_�@Diag S?ummary<_IJ�
CONSLOG�1__&Q_�_NQC�onsole l�og�_HK	TPA'CCN�_o%o?o�JUTP Acc?ountin�_IJ�FR6:IPKDMP.ZIPso�wH
�o�oKU[`Exception�o�yk'PMEMCHECCK5o�_*_K�Q�Memory D�ataL�F!l{�)6qRIPE�_p$6�Zs%�q� Packet yL�_�DL�$�	r�qSTAT����S� %�rS�tatusT��	FTP���:���Vw��Qmment �TBD؏� >I�)ETHERN�E���
q�[�NQ?Ethern�p�P?figura�oOD~DCSVRF̏в�ďݟd��� v�erify al�l��{D}.���DIFF՟��͟b��s��diffd��
q>��CHG01Y�@��R��f�z���-?��2ݯį֯k�v������3a�H�Z��� ��ϥ�VT�RNDIAG.LAS�̿޿s�^q3�O Ope���q SQ�nosticEW0��)VDEV7�DATt�Q�c�u��g�Vis��De�vice�Ϫ�IM�G7ºo����y��s��Imagߨ��UP��ES��T��FRS:\�� ��OQUpdates� List �IJ�g�FLEXEVEANQ�X�j߃�f�F� UIF Ev����B,�s�)
�PSRBWLD.CM��sL�������PPS_ROBO�WEL��GLo�G�RAPHICS4�Dy�b�t��%�4D Graph�ics File�u��AOɿ�rG�IG���u�
Yv�GigE�ة�BNߵ? )��HADOW�����\s�Shadow �Chang���v�bQRCMERAR�n�\s� �CFG Erro�r�tail� �MA��CMSGLIB���"^o� ��T7�)�ZD�����/XwZD6 a�d�HPNOT�I���
/�/ZuN?otific��H/��AGUO�/yO? �O'?P?OOt??�?�? 9?�?]?�?O�?(O�? LO^O�?�OO�O5O�O �OkO _�O$_6_�OZ_ �O~_�__�_C_�_�_ y_o�_2o�_?oho�_ �oo�o�oQo�ouo
 �o@�odv� )�M����� <�N��r������7� ̏[������&���J� ُW������3�ȟڟ i�����"�4�ßX�� |������A�֯e�� ���0���T�f����� �����O��s��� ��>�Ϳb��oϘ�'� ��K����ρ�ߥ�:� L���p��ϔߦ�5��� Y���}���$��H��� l�~���1�����g� ��� �2���V���z� 	�����?���c���
 ��.��Rd��� ��M�q� <�`���%� I��/�8/J/ �n/��/!/�/�/W/ �/{/?"?�/F?�/j?�|??�?/?�?�?�$�FILE_FRS�PRT  ����0�����8MDONLY� 1]�5�0 �
 �)MD:�_VDAEXTP.ZZZ�?�?_OnK�6%NO �Back fil�e 9O�4S�6P e?�OOO�O�?�O__? >_�Ob_t__�_'_�_ �_]_�_�_o(o�_Lo �_po�_}o�o5o�oYo �o �o$�oHZ�o ~��C�g� �	�2��V��z��� ���?�ԏ�u�
����.�@��4VISBC�KHA&C*.V�DA�����FR:�\Z�ION\DA�TA\v�����Vision VD�B��ŏ���'�5� �Y��j������B� ׯ�x����1���ү g�������X���P�� t���Ϫ�?�οc�u� ϙ�(Ͻ�L�^��ς� �)���M���q� ߂� ��6���Z�����%����I�������:LU�I_CONFIG7 ^�5m��� $ h�F{ �5������)�;�I���|xq�s������� ����a��� $6 ��Gl~���K ��� 2�V hz���G�� �
//./�R/d/v/ �/�/�/C/�/�/�/? ?*?�/N?`?r?�?�? �???�?�?�?OO&O �?JO\OnO�O�O)O�O �O�O�O�O_�O4_F_ X_j_|_�_%_�_�_�_ �_�_o�_0oBoTofo xo�o!o�o�o�o�o�o �o,>Pbt� ������� (�:�L�^�p������ ��ʏ܏���$�6� H�Z�l��������Ɵ ؟ꟁ�� �2�D�V� h���������¯ԯ� }�
��.�@�R�d��� ��������п�y�� �*�<�N�`����ϖ� �Ϻ�����u���&� 8�J���[߀ߒߤ߶� ��_������"�4�F� ��j�|������[� ������0�B���f� x���������W����� ,>��bt� ���O���(:�  x�FS�$FLUI�_DATA _�������uRESU_LT 2`��� �T�/�wizard/g�uided/st�eps/Expertb��//+/�=/O/a/s/�/�/�*��Continu�e with G�ance�/�/�/ ??(?:?L?^?p?�?,�?�? T-U�>�90 �� �?؅��9��ps �?0OBOTOfOxO�O�O �O�O�O�O�O� �_ /_A_S_e_w_�_�_�_ �_�_�_�_n�?�?�?:�<Frip�O o�o�o�o�o�o�o�o !3E_i{� �������� /�A�S�o$on�HoA�O�TimeUS/DST[���� ��+�=�O�a�s�������'Enabl �/˟ݟ���%�7�@I�[�m������T��?{�ݯ����Æ24Ώ3�E�W�i�{��� ����ÿտ翦���� /�A�S�e�wωϛϭ� �������ϴ�Ưد�� G��Region�χߙ߽߫����������)�;�+A?mericasou� ������������ �)�;��?�y�#����G�Y��ditorL�������#5�GYk}��+ T�ouch Pan�el �� (re�commen�) ���*<N `r��U��e�w���������accesd�./@/R/d/v/�/��/�/�/�/�/Q|C�onnect t�o Network�/(?:?L?^?p?�?��?�?�?�?�?�?Y��B������!/���Introducts߆O�O�O�O�O �O�O__(_:_U^_ p_�_�_�_�_�_�_�_` oo$o6oHo e� Oeo?O�X_�o�o�o �o'9K]o ��R_����� �#�5�G�Y�k�}���"��h`�ooj}oߏ �o��*�<�N�`�r� ��������̟ޟ�� �&�8�J�\�n����� ����ȯگ쯫���Ϗ 1��X�j�|������� Ŀֿ�����0�� A�f�xϊϜϮ����� ������,�>���_� !���E��߼������� ��(�:�L�^�p�� ��߸������� �� $�6�H�Z�l�~���O� ��s������� 2 DVhz���� ����
.@R dv������ ��/��'/���`/r/ �/�/�/�/�/�/�/? ?&?8?�\?n?�?�? �?�?�?�?�?�?O"O 4O�UO/yO�OO?�O �O�O�O�O__0_B_ T_f_x_�_I?�_�_�_ �_�_oo,o>oPobo to�oEO�OiO�o�o�O (:L^p� ������_ �� $�6�H�Z�l�~����� ��Ə؏�o�o�o�/� �oV�h�z������� ԟ���
��.��R� d�v���������Я� ����*������ ��C�����̿޿�� �&�8�J�\�nπ�?� �϶����������"� 4�F�X�j�|ߎ�M�_� q��ߕ�����0�B� T�f�x�������� ������,�>�P�b� t��������������� ����%��L^p� ������  $��5Zl~�� �����/ /2/ ��S/w/9�/�/�/ �/�/�/
??.?@?R? d?v?�?�/�?�?�?�? �?OO*O<ONO`OrO �OC/�Og/�O�/�O_ _&_8_J_\_n_�_�_ �_�_�_�_�?�_o"o 4oFoXojo|o�o�o�o �o�o�O�o�O�O�o Tfx����� ����,��_P�b� t���������Ώ��� ��(��oI�m�� C�����ʟܟ� �� $�6�H�Z�l�~�=��� ��Ưد���� �2� D�V�h�z�9���]��� ѿ����
��.�@�R� d�vψϚϬϾ��Ϗ� ����*�<�N�`�r� �ߖߨߺ��ߋ�տ�� ��#��J�\�n��� ������������"� ��F�X�j�|������� ������������ ��u7���� ��,>Pb t3������� //(/:/L/^/p/�/ ASe�/��/ ?? $?6?H?Z?l?~?�?�? �?�?��?�?O O2O DOVOhOzO�O�O�O�O �O�/�/�/_�/@_R_ d_v_�_�_�_�_�_�_ �_oo�?)oNo`oro �o�o�o�o�o�o�o &�OG	_k-_� �������"� 4�F�X�j�|������ ď֏�����0�B� T�f�x�7��[�� �����,�>�P�b� t���������ί��� ��(�:�L�^�p��� ������ʿ��뿭�� џӿH�Z�l�~ϐϢ� ����������� �߯ D�V�h�zߌߞ߰��� ������
��ۿ=��� a�s�7ߚ������� ����*�<�N�`�r� 1ߖ����������� &8J\n-�w� Q������" 4FXj|��� �����//0/B/ T/f/x/�/�/�/�/ ���/?�>?P?b? t?�?�?�?�?�?�?�? OO�:OLO^OpO�O �O�O�O�O�O�O __ �/�/�/?i_+?�_�_ �_�_�_�_�_o o2o DoVoho'O�o�o�o�o �o�o�o
.@R dv5_G_Y_�}_� ���*�<�N�`�r� ��������yoޏ��� �&�8�J�\�n����� ����ȟ����� 4�F�X�j�|������� į֯����ˏ�B� T�f�x���������ҿ �����ٟ;���_� !��ϘϪϼ������� ��(�:�L�^�p߁� �ߦ߸������� �� $�6�H�Z�l�+ύ�O� ��s�������� �2� D�V�h�z��������� ������
.@R dv����}�� �����<N`r �������/ /��8/J/\/n/�/�/ �/�/�/�/�/�/?� 1?�U?g?+/�?�?�? �?�?�?�?OO0OBO TOfO%/�O�O�O�O�O �O�O__,_>_P_b_ !?k?E?�_�_{?�_�_ oo(o:oLo^opo�o �o�o�owO�o�o  $6HZl~�� �s_�_�_���_2� D�V�h�z������� ԏ���
��o.�@�R� d�v���������П� �������]�� ��������̯ޯ�� �&�8�J�\������ ����ȿڿ����"� 4�F�X�j�)�;�M��� q���������0�B� T�f�xߊߜ߮�m��� ������,�>�P�b� t�����{ύϟ� ���(�:�L�^�p��� ������������ �� 6HZl~�� �������/ ��S�z���� ���
//./@/R/ d/u�/�/�/�/�/�/ �/??*?<?N?`? �?C�?g�?�?�?O O&O8OJO\OnO�O�O �O�Ou/�O�O�O_"_ 4_F_X_j_|_�_�_�_ q?�_�?�_�?�_0oBo Tofoxo�o�o�o�o�o �o�o�O,>Pb t������� ��_%��_I�[��� ������ʏ܏� �� $�6�H�Z�~����� ��Ɵ؟���� �2� D�V��_�9�����o� ԯ���
��.�@�R� d�v�������k�п� ����*�<�N�`�r� �ϖϨ�g��������� ��&�8�J�\�n߀ߒ� �߶��������߽�"� 4�F�X�j�|���� ��������������� Q��x����������� ����,>P� t������� (:L^�/� A��e���� // $/6/H/Z/l/~/�/�/ a�/�/�/�/? ?2? D?V?h?z?�?�?�?o ���?�O.O@ORO dOvO�O�O�O�O�O�O �O�/_*_<_N_`_r_ �_�_�_�_�_�_�_o �?#o�?Go	Ono�o�o �o�o�o�o�o�o" 4FXio|��� ������0�B� T�ou�7o��[o��ҏ �����,�>�P�b� t�������iΟ��� ��(�:�L�^�p��� ����e�ǯ��믭��� $�6�H�Z�l�~����� ��ƿؿ����� �2� D�V�h�zόϞϰ��� �����Ϸ��ۯ=�O� �v߈ߚ߬߾����� ����*�<�N��r� ������������ �&�8�J�	�S�-�w� ��c���������" 4FXj|��_� ����0B Tfx��[���� ����/,/>/P/b/ t/�/�/�/�/�/�/�/ �?(?:?L?^?p?�? �?�?�?�?�?�?�� ��EO/lO~O�O�O �O�O�O�O�O_ _2_ D_?h_z_�_�_�_�_ �_�_�_
oo.o@oRo O#O5O�oYO�o�o�o �o*<N`r ��U_����� �&�8�J�\�n����� ��couo�o鏫o�"� 4�F�X�j�|������� ğ֟蟧���0�B� T�f�x���������ү ������ُ;���b� t���������ο�� ��(�:�L�]�pς� �Ϧϸ������� �� $�6�H��i�+���O� ����������� �2� D�V�h�z���]��� ������
��.�@�R� d�v�����Y߻�}��� �ߣ�*<N`r ��������� &8J\n�� �������/�� 1/C/j/|/�/�/�/ �/�/�/�/??0?B? f?x?�?�?�?�?�? �?�?OO,O>O�G/ !/kO�OW/�O�O�O�O __(_:_L_^_p_�_ �_S?�_�_�_�_ oo $o6oHoZolo~o�oOO �OsO�o�o�O 2 DVhz���� ���_
��.�@�R� d�v���������Џ� �o�o�o�o9��o`�r� ��������̟ޟ�� �&�8��\�n����� ����ȯگ����"� 4�F���)���M��� Ŀֿ�����0�B� T�f�xϊ�I������� ������,�>�P�b� t߆ߘ�W�i�{��ߟ� ��(�:�L�^�p�� ������������ $�6�H�Z�l�~����� ������������/ ��Vhz���� ���
.@Q dv������ �//*/</��]/ �/C�/�/�/�/�/? ?&?8?J?\?n?�?�? Q�?�?�?�?�?O"O 4OFOXOjO|O�OM/�O q/�O�/�O__0_B_ T_f_x_�_�_�_�_�_ �_�?oo,o>oPobo to�o�o�o�o�o�o�O �O%7�_^p� ������ �� $�6��_Z�l�~����� ��Ə؏���� �2� �o;_���K�� ԟ���
��.�@�R� d�v���G�����Я� ����*�<�N�`�r� ��C���g���ۿ��� �&�8�J�\�nπϒ� �϶����ϙ����"� 4�F�X�j�|ߎߠ߲� ���ߕ�����˿-�� T�f�x�������� ������,���P�b� t��������������� (:���� A�����  $6HZl~=�� �����/ /2/ D/V/h/z/�/K]o �/��/
??.?@?R? d?v?�?�?�?�?�?� �?OO*O<ONO`OrO �O�O�O�O�O�O�/�O �/#_�/J_\_n_�_�_ �_�_�_�_�_�_o"o 4oE_Xojo|o�o�o�o �o�o�o�o0�O Q_u7_���� ����,�>�P�b� t���Eo����Ώ��� ��(�:�L�^�p��� A��eǟ��� �� $�6�H�Z�l�~����� ��Ưد����� �2� D�V�h�z�������¿ Կ�������+��R� d�vψϚϬϾ����� ����*��N�`�r� �ߖߨߺ�������� �&��/�	�S�}�?� ������������"� 4�F�X�j�|�;ߠ��� ��������0B Tfx7��[�� ���,>Pb t�������� //(/:/L/^/p/�/ �/�/�/�/���� !?�H?Z?l?~?�?�? �?�?�?�?�?O O� DOVOhOzO�O�O�O�O �O�O�O
__._�/�/ ?s_5?�_�_�_�_�_ �_oo*o<oNo`oro 1O�o�o�o�o�o�o &8J\n�?_ Q_c_��_���"� 4�F�X�j�|������� ď�oՏ����0�B� T�f�x���������ҟ ����>�P�b� t���������ί�� ��(�9�L�^�p��� ������ʿܿ� �� $��E��i�+��Ϣ� ����������� �2� D�V�h�z�9��߰��� ������
��.�@�R� d�v�5ϗ�Yϻ�}�� ����*�<�N�`�r� �������������� &8J\n�� �������� ��FXj|��� ����//��B/ T/f/x/�/�/�/�/�/ �/�/??�#�G? q?3�?�?�?�?�?�? OO(O:OLO^OpO// �O�O�O�O�O�O __ $_6_H_Z_l_+?u?O? �_�_�?�_�_o o2o DoVohozo�o�o�o�o �O�o�o
.@R dv����}_�_ �_�_��_<�N�`�r� ��������̏ޏ��� ��o8�J�\�n����� ����ȟڟ����"� ���g�)������� į֯�����0�B� T�f�%���������ҿ �����,�>�P�b� t�3�E�W���{����� ��(�:�L�^�p߂� �ߦ߸�w����� �� $�6�H�Z�l�~��� �����������2� D�V�h�z��������� ������
-�@R dv������ ���9��]� �������/ /&/8/J/\/n/-�/ �/�/�/�/�/�/?"? 4?F?X?j?)�?M�? qs?�?�?OO0OBO TOfOxO�O�O�O�O/ �O�O__,_>_P_b_ t_�_�_�_�_{?�_�? oo�O:oLo^opo�o �o�o�o�o�o�o  �O6HZl~�� �������_o �_;�e�'o������ ԏ���
��.�@�R� d�#��������П� ����*�<�N�`�� i�C�����y�ޯ�� �&�8�J�\�n����� ����u�ڿ����"� 4�F�X�j�|ώϠϲ� q�������	�˯0�B� T�f�xߊߜ߮����� �����ǿ,�>�P�b� t����������� ��������[�߂� ������������  $6HZ�~�� ����� 2 DVh'�9�K��o� ���
//./@/R/ d/v/�/�/�/k�/�/ �/??*?<?N?`?r? �?�?�?�?y�?��? �&O8OJO\OnO�O�O �O�O�O�O�O�O_!O 4_F_X_j_|_�_�_�_ �_�_�_�_o�?-o�? QoOxo�o�o�o�o�o �o�o,>Pb !_������� ��(�:�L�^�o� Ao��eog�܏� �� $�6�H�Z�l�~����� ��s؟���� �2� D�V�h�z�������o� ѯ�����˟.�@�R� d�v���������п� ���ş*�<�N�`�r� �ϖϨϺ�������� ����/�Y���ߒ� �߶����������"� 4�F�X��|���� ����������0�B� T��]�7߁���m��� ����,>Pb t���i���� (:L^p� ��e�w�������� $/6/H/Z/l/~/�/�/ �/�/�/�/�/� ?2? D?V?h?z?�?�?�?�? �?�?�?
O���OO /vO�O�O�O�O�O�O �O__*_<_N_?r_ �_�_�_�_�_�_�_o o&o8oJo\oO-O?O �ocO�o�o�o�o" 4FXj|��__ ������0�B� T�f�x�������moϏ �o�o�,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� ��� !��E��l�~����� ��ƿؿ���� �2� D�V��zόϞϰ��� ������
��.�@�R� �s�5���Y�[����� ����*�<�N�`�r� ����g�������� �&�8�J�\�n����� ��c�����������" 4FXj|��� ������0B Tfx����� ��������#/M/ t/�/�/�/�/�/�/�/ ??(?:?L?p?�? �?�?�?�?�?�? OO $O6OHO/Q/+/uO�O a/�O�O�O�O_ _2_ D_V_h_z_�_�_]?�_ �_�_�_
oo.o@oRo dovo�o�oYOkO}O�O �o�O*<N`r ��������_ �&�8�J�\�n����� ����ȏڏ����o�o �oC�j�|������� ğ֟�����0�B� �f�x���������ү �����,�>�P���!�3������$FM�R2_GRP 1�a��� ��C4  B]�[�	 [�߿��ܰE�� F;@ 5W�S��ܰJ��NJk��I'PKHu���IP�sF!�=��?�  W�S��ܰ9�<9���896C'�6<,5��=�A�  �Ϲ�BHٳB�հ�����@�33�33�S�۴��ܰ@UUT'�@��8��W��>u.�>*���<����=[��B=���=|�	<�K�<�q߼=�mo����8�x	7H�<8�^6�Hc7��x?���� ������"��F�X���_CFG b»T Q����X�NO º�
F0�� ��W�R�M_CHKTYP  ��[�ʰ̰��ROM�_MI�N�[���9�����X��SSBh�c��� �ݶf�[�]����^�TP_DEF_O��[�ʳ��IRC�OM���$GE�NOVRD_DOr.�d���THR.�� dd��_EN�B�� ��RAV�C��dO�Z� ����Fs  G!�� GɃ�I��C�I(i J�C��+���%������ �QOU*��j¼������<6�i�C��;]�[�C�  �D�+��@���B����.\��R SMT��k_	�ΰ\��$HOS�TCh�1l¹[�s�d�۰ MC[����/Z� _ 27.0� 1�/  e�/??'? 9?G:�/j?|?�?�?�,�Z?T3	anonymouy �?�?	OO -O?N�/ڰRHRK�/ �?�O�/�O�O�O�O_ V?3_E_W_i_�O&_�? �_�_�_�_�_@O�_dO vOSo�_�Ojo�o�o�o �o_�o+=`o �_�_�����o &o8oJoL9��o]�o� �������oɏۏ��� �4�j+�Y�k�}��� ������ ��T� 1�C�U�g��������� ��ӯ��x�>��-�?� Q�c�����Ο���Ͽ ����)�;ς�_� qσϕϧ�ʿ ���� ��%�7�~������ �ϣ������������ ��3�E�W�i�ߍ��� ����������@�R�d� v�x�J��߉������� �����+=`� �������:$~h!ENT 1m� P!V  7 ?.c& �J�n���/ �)/�M//q/4/�/ X/j/�/�/�/�/?�/ 7?�/?m?0?�?T?�? x?�?�?�?O�?3O�? WOO{O>O�ObO�O�O �O�O�O_�OA__e_ (_:_�_^_�_�_�_�ZQUICC0�_�_�_?od1@oo.o��od2�olo~o�o!ROUTER�o��o�o/!PCJ�OG0!1�92.168.0�.10	o�SCAMgPRT�\!pu11yp��vRT�o���� !Sof�tware Op�erator Panel�mn��NAME !�
?!ROBO�v��S_CFG 1l��	 ��Auto-sta�rted'�FTP2��I�K2�� V�h�z�������ԟ ����	���@�R�d� v���	������� :���)�;�M�_�&��� ������˿�p��� %�7�I�[��"�4�F� ڿ��������!�3� ��W�i�{ߍߟ���D� ��������/�vψ� ��w�ߛ��Ͽ����� ����+�=�O�a��� �������������8� J�\�n�p�]��� �������# 5X�k}��� �0/D1/x U/g/y/�/RH/�/�/ �/�//?�/??Q?c? u?�?���/?�? :/O)O;OMO_O&?�O �O�O�O�O�?pO__ %_7_I_[_�?�?�?t_ �O�_O�_�_o!o3o �OWoio{o�o�_�oDo��o�o�o����_?ERR n��-�=vPDUSIZ � �`^�P�Tt�>muWRD ?�΅�Q�  ?guest�f�������~�SC�DMNGRP 2�o΅Wp���Q�`���fKL� �	P01.05� 8�Q   ��|��  ;�|��  z[ ����w���*����Ť�x����[ݏȏ��+בPԠ�������)����D�r����؊p"�PlJ�P���Dx��dx��*�����%�_GROUU7�pLyN��q	/�o���QUP���UTu� �TY�àL}?pTTP�_AUTH 1q�L{ <!iP�endan�����o֢!KARE�L:*������K�C��ɯۯ��VI�SION SET �9����P�>�h�� f����������ҿ�����X�CTRL� rL}O�uſa
��aFFF9E�3-ϝTFRS:DEFAULT���FANUC �Web Server�ʅ�u�X���t @���1�C�U�g�;t�WR_CONFI�G s;� ���=qIDL_CP�U_PC���aB�ȠP�� BH��M�IN�܅q��GNR_IOFq{r�`Rx���NPT_SIM_�DO��STA�L_SCRN� ��.�INTPMODNTOLQ����RTY0����-�\��ENBQ�-���O�LNK 1tL{ �p������)�;�M�>��MASTE�%����SLAVE �uL|�RAMCA�CHEk�c�O^�O�_CFG������U�OC�����CMT_�OP���PzYC�L������_ASG� 1v;��q
  O�r������ �&8J\W��ENUMzsPy
���IP����RTRY_CN��M�=�zs���Tu ������w���p/�p��P�_MEMBERSg 2x;�l� $��X"��?�Q'W/i)���RCA_ACC� 2y�  X�cN �e��b'63`�"��Q�&�#�#�/�!�/c�!�BUF001 2�z�= cu0  u0c+:4�;:4N:4XF� � F�^�:3^�V:3_j4j4%j4U6j4Hj4Xj4jj4}z:3` � �0�`�4"�42�4D��4T�4g�4w�4���4��4��4��4�j�4�4�:3a"DY"D�4a5"DG"DeW"Di"D�4a�"DU�"D�"D�"D�"D��"D�:3b�D��D'�D8�DJ�DZ��Dl�D}�D��D���D��DĚDԚD�J�D�:4	:392$? 63:1@1ERI0ERQ0ER Y0Z1`1:1h1:1p1uR y0uR�0uR�0uR�0uR �0uR�0uR�0:1�1�1 �1�R�0�R�0�R�0�R �0�R�0�R�0�R�0�R �0�R@�R	@�R@�R @�R!@:1(A-b1@-b �T@A-bI@-bQ@-bY@ -b�ThA-bq@-by@-b �@-b�@-b�@-b�@:1 �A�b�@�b�@�b�@�b �@�b�@�b�@�b�@�b �@�b�@�b�@�b�@�b P�b	P�bPERP:193-_65GSNrI2WS NrY2gSnri2wS~ry2 �S~r�2�S~r�2�S~r �2�S�r�2�S�r�2�S �r�2�S�r�2�S�r�2 c�r	Bc�rB'c�� (C7c6��t@COc6�QB _c6��thCwc6�yB�c 6��B�c6��B�c���B �c���B�c���B�c�� �B�c���B�c���Bs���	RsNrR'v��2E{�4r�}ŋ����<����o�o��2�H�IS!2}� ���! 2024-O06-1O������П���  �� �9 X��o��";�WQ�(�:�L�^�o�X7�mv��06�������Ư�����Z؞M 9 hL!��mv��;M ��1�C� r�O�!���������� ο����(�_�q� ^�pςϔϦϸ����� �� �7�I�6�H�Z�l� ~ߐߢߴ������!� � �2�D�V�h�z�� ����������
�� .�@�R�d�v���k�� ,P������������U:�b�:��a� &�d� A_q��q���������&�  @�A��;��c��b�o�c �CUg����t� ����	//-/?/ v���/�/�/�/�/ �/�/??)?`/r/_? q?�?�?�?�?�?�?�? O8?J?7OIO[OmOO �O�O�O�O�OO"O_ !_3_E_W_i_{_�_�_ �_����5p�����o�$o6o���B��B� ^secro�o�o�o�� o�oݪXc�b��"k� ��Br�d v��O�O�o��� ��*�<�N�`�r�� �����̏ޏ���� &�8�J����������� ��ȟڟ����"�Y� k�X�j�|�������į ֯���1�C�U�B�T� f�x���������ҿ�_���I_CFG 2�~�[ H
C�ycle Tim}e�Busy��Idl��m�in�S�U�p��Read>(�DowG�C��: X��Coun}t�	Num �"������`����oPROG���U��P�)/so�ftpart/g�enlink?c�urrent=m�enupage,?1133,1�C��U�g�y�Tä�SDT�_ISOLC  ��Y� ���J�23_DSP_ENB  ��T���?INC ����c���A   ?� � =���<#��
���:�o ��2�D��a/�l���OB��C��O��ֆ��G_GROUP �1���-d<�*�����t�?"�����`Q'�L� ^�p�/�����������\�~�G_IN_�AUTO����PO�SRE���KANJI_MASK0���DRELMONG ��[���by�� ������f��%������d-���KCL_L N�UM��G$KEYLOGGINGD��P�������LAN�GUAGE ��U��DE?FAULT ��Q�LG�����S�U��ax�Hp8T�oH  ��`'0����`;�`JrK��e;���
*!(UTg1:\ J/ L/ Y/k/}/�/�/�/�/�/��/�/$>(�H?�VL�N_DISP ����P�&�$�^4OCgTOL�0�aDz�����
�1GBOOK ��d4V�11�07u%O!O3O EOWOiKyM�TËIgF	�5)����O}����2_BUFF ;2��� ��`2O�_�2��6_M�R_ d_�_�_�_�_�_�_�_ �_o3o*o<oNo`o�o��o�o�o���ADCS ������L�O���+=Oa�dI�O 2��k +������� �����*�:�L� ^�r���������ʏ܏����$�6�J�uuE_R_ITM��d�� ����ǟٟ����!� 3�E�W�i�{��������ïկ�����7x�S�EVD��t�TYP����s�������)RSTe�eSC�RN_FL 2�
�}�����/�`A�S�e�wϨ�TP{���b��=NGNA�M��E��dUPS�f0GI��2�����_LOAD��G� %��%PI�CKUP_PRE�NSA�Ϭ6MAXUALRMb2�@���
K���+��Ģ2  �3�AK�Ci0���qO=_'X�Ӭ�Pw 2��; �*V�	����
* � ��4��*��'�`�	x N��z�������� ���1�C�&�g�R��� n�����������	 ��?*cFX�� �����; 0q\���� ���/�/I/4/ m/X/�/�/�/�/�/�/ �/�/!??E?0?i?{? ^?�?�?�?�?�?�?�? OOAOSO6OwObO�O�D�DBGDEF ���գѢѤO�@_LDXDISA�����ssMEMO_A�P��E ?��
 �A�H$_6_H_�Z_l_~_�_�_K�FR�Q_CFG �ږ��CA �G@�4�S�@<��d%�\o�_�P�Ґ��^��*Z`/\b **:eb�DXojh o�F�o�o�o�o�o �o;�O��dZ�U0�y|��z,(9� Mt���1��B�g� N���r��������̏�	���?�A�ISCg 1���K` ��O �����O���O֟�����K�]�_MSTR ��3��SCD 1�]��l�� {�����دïկ��� 2��V�A�z�e����� ��Կ�������@� +�=�v�aϚυϾϩ� ��������<�'�`� K߄�oߨߓߥ����� ���&��J�5�Z�� k����������� ���F�1�j�U���y� ������������0`T?x�MK�Q��,��Q�$MLoTARM�R�?g� ~s�@�|��@METPU�@�l��4�NDSP_ADCOL��@!CMNT7 �*FNSW(F�STLIxi%� �,����Q���*POSCF��bPRPMV�S�T51�,� 4�R#�
g!|qg%w/ �'c/�/�/�/�/�/�/ ?�/?G?)?;?}?_?�q?�?�?�?�?�1*S�ING_CHK � {$MODA��S�e���#ED�EV 	�J	�MC:WLHSIZ�E�Ml �#ETAS�K %�J%$1�23456789� �O�E!GTRIGw 1�,� l�E�o#_�y_S_�}�FY�P�A�u9D"CEM_INF 1�?k�`)AT&�FV0E0X_�])��QE0V1&A�3&B1&D2&�S0&C1S0=>�])ATZ�_#o
dH'oOo�QC_wohAo�obo�o�o�o �_&�_�_�_o� 3o��o���o�� "�4��X���A Se֏���C�0� ��f�!���q����� s�䟗�����͏>�� b���s���K���w�� �ٯ�ɟ۟L���� #�����Y�ʿ�� ��$�߿H�/�l�~�1� ��U�g�y����ϯ� � 2�i�V�	�z�5ߋ߰������PONITOR�G ?kK   �	EXEC1To�2�3�4�Q5��@�7�8�9o���� (��4��@��L�� X��d��p��|��U2��2��2��2��U2��2��2��2��U2��2��3��3���3(�#AR_GRP�_SV 1��[� (�1���?��C�=@�H���! ?gc�"RM�A_Ds���N��ION_DB�-@�1Ml  ��� �� �JD"�� �/�  ��FH��N   ,��c �/�FI-ud1}E���)�PL_NAME �!�E� �!�Default �Personal�ity (fro�m FD)b (R�R2�� 1�L?�XL�p�X  d�-?Q cu������ �//)/;/M/_/q/�/�/�/EC2)�/�/ �/??,?>?P?b?t?EB<�/�?�?�?�?�? �?
OO.O@OROdO�%�6�?�N
�O�O�P�O�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_�O�O2oDoVo hozo�o�o�o�o�o�o �o
.@o!ov �������� �*�<�N�`�r������ Fs  GT�G�M���  �ÏՍ�d�������(�6� �����
 �m�~�h����� ������ğ ֟�����:���
�]�4m����	`�������į��:�oA������ A�  /���P��� �r�������^�˿ݿ�ȿ��%��R�� �1��	X ��, � ��� a�g @Dj t�?�z��`�?� |��A/���t�{	��;�	l���	 �xoJ����� �� �<�@����� ��·�K��K ��K=�*�J���J�?��J9���
�ԏC߷�@�t��@{S�\��(E�hє��.��I���ڌ���T�;f�ґ�$��3���´  �@���>�Թ�$�  >̿���ӧU��g�x`���� ��
���Ǌ��� ��  {  �@T�����  ��O �l�ϊ�-�	�'� � ���I� �  y�<�+�:�È��?È=�����0����N �[��n @���f����f�k���,�av� � '��Yэ�@2��@�0@�Ь����C��Cb C���\C�������G�@�� %! ����� )�Bb $/�!��L�Dz�o�ߓ~���0��( �� -��������!9�D� � 9�恀?�fafG�*<� }��q�1�89��>���bp��(�(9��P���	������>�?���9�x9�W�<�
6b<߈;�܍�<�ê<���<�^��dI/��A�{��f�|��,�?fff?_��?&� T�@�.��"�J<?�\��"N\�6���!�� (�|��/z��/j'��[ 0??T???x?c?�?�?��?�?�?�?6��%F ���?2O�?VO�/wO�)�IO�OEHG@ G�@09�G�� G}ଙO�O�O_	_B_�-_f_Q_BL9�B��Aw_[_�_b��_�[ �_��mO3o�OZo�_~o�o�o�o���b��PV( @|po	lo@-*cU�ߡA���r59�CP�Lo�}?����#�l�6��W9���6�3Cv�q�CH3� jD�t����q�����|^�(hA� �A�LffA]��??�$�?��;��°u�æ�)��	ff��Cϼ#�
���g\�)�"�33C�
������<����؎G�B����L�B�s����	"�;�H�ۚG���!G��WIY�E���C�+��8�I۪I��5�HgMG��3E��RC��j=x�
�pI����G��fIV�=�E<YD �C<�ݟȟ����7� "�[�F��j������� ٯį���!��E�0� i�T�f�����ÿ��� ҿ����A�,�e�P� ��tϭϘ��ϼ���� ��+��O�:�s�^߃� �ߔ��߸������ � 9�$�6�o�Z��~�� �����������5� � Y�D�}�h����������������
C.(�䁳��/"��<�<��t��q3�8����q�4Mgu���q��VwQ�
4p�+4�]$$d@R�v���uPD"	P��Q�_/Z/0=/(/a/L+Rg/n/`�/�/�/�/�/  %��/�/+??O?:?s?�/�_�?�?�?�; �?�?O�? OFO4O�rLO^O�O�O�O�O�O��J  2 FsޙwGT�V��M�uBO�|r�pp�C��S@�R_�poy_��_^_�_o \!�WɃ�_oo(o~�z?���@@�z��D�p�pk1:�p�~
 6o�o �o�o�o�o�o)�;M_q�ڊsa �����D���$MR_CABL�E 2�� S]��T�La�Ma?�PMaLb�p��Z��&P�C�p?aO4>�B���?b�w	$?`?aE��F�?f��v�l � ��&P�v�wdN��{0��$��n?`�F:�H( 6�H�XT��6P?`�C!��Č���n�ə�&�ˡ(͂���| ��&P���C���=�����n�
9��z��� �bڅ��s9��T�,� >���b�������Ɵ�� Ο3�.��P�(�:��� ^���j��#?`���� ��<h�H�Z�l�<hw*��** �s�OM ��y����B?b�$%�% 234567O8901ɿ۵ ƿH���?`�?`AQ?`�?a
�z�n�ot sent 앺�W�T�ESTFECSA�LG� eg;jAQdȎ�ga%�
���@��?d�r�̹�������� 9UD1:�\mainten�ances.xm�S�.�@�vj�DEFAULT�\~�rGRP 2����  phd�G?e � �%1st �mechanic�al checkl�?a���������E��Z�(�:��L�^�?b��cont?roller�Ԍ��߰��D����� ��$�s�M��L�?b�"8b���v��B������������/�C }�a�6����d�v���s�C��g�e��. batt�ery�&��E	 S(:L^p�	|��duiz�ablet  D�а!�!���D��/"/�4/s��greaYs�>gf�r#-?`|!�/�E��/�/�/h�/�/s�
�oi,�g/y/�/�/t?�?�?�?�?s��
�?f	�W��1<?`AO�E
c?8OJO\OnO�O�!t��?O��'O�O�_ _2_D_s�Ov�erhauE��L��R x?`�Q�_���O�_�_�_�_o?`A$�_0o����_o �_ �o�o�o�o�oo�o?o QocoJ\n�� �o�)��"� 4�F���|��k�� ď֏����[�0�B� ��f�����������ҟ !���E�W�,�{�P�b� t�����矼���� A��(�:�L�^����� ѯ㯸��ܿ� �� $�s�Hϗ���~�Ϳ�� ��������9��]�o� Dߓ�h�zߌߞ߰��� ��#�5�G���.�@�R� d�v��ߚ�������� ����*�y���`��� O������������?� &u�J��n�� ���);_ 4FXj|��� �%�//0/B/ �f/���/��/�/ �/�/?W/,?{/�/b? �/�?�?�?�?�??�? A?S?(Ow?LO^OpO�O �O�?�OOO+O�O_ $_6_H_Z_�O~_�O�O �O�_�_�_�_o o�PeR	 T"oOoaoso �_�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z��������ԏ���
�� � ��Q?�  @eQ �oW�i�{��eVC�����̟bX*�** �Q�V�� � �2�D��h�z��������_�S��� ���կ7�I�[��� ��ɯ/���ǿٿ#�� �!�3�}�����{ύ� ���s�������C�U� g��S�e�w�9ߛ߭�п�	��eUeQ�$�MR_HIST �2��U�� 
� \jR$ 2345678901*�(2����)�9c_�� ��R��a_������� ��=�O�a��*�x��� ��r�������9 ��]o&�J�� ���#�G��k}4�Z�SK�CFMAP  .�U�����Z��ONR�EL  �����лEXCFE�NB'
��!F�NC$/$JOGO/VLIM'd�m ��KEY'p%y%_PAN(�"�"��RUN`,p%��SFSPDTY�PD(%�SIGN|/$T1MOTb/�!�_CE_G�RP 1��U �"�:`��n?Z[?�? �؆?�?~?�?�?�?!O �?EO�?:O{O2O�O�O hO�O�O�O_�O/_�O (_e__�_�_�_�_v_��_�_�_o�׻QZ_EDIT4��#�TCOM_CFG 1��'%to�o��o 
Ua_ARC�_!"��O)T_M�N_MODE6=�Lj_SPL�o2&UAP_CPL�o�3$NOCHECK� ?� � Rdv��� ������*�<��N�`��NO_WA�IT_L 7Jg50N�T]a���UZ޲�_ERR?12���ф��	��-�����R�d����`O�����| �f
a�����A����/^$C3������BL��<� �� ?�j�ϟj�����قPARAM�Ⴓ��N��
oQ�h�o��� = e������گ� ȯ��"�4��X�j�F�g蜿��A�ҿ�"?ODRDSP�c6�/(OFFSET_�CAR@`�o�DI�S��S_A�`A�RK7KiOPEN_FILE4�1�a�Kf�`OPTION�_IO�/�!��M_�PRG %�%c$*����h�WOT�[�E7O��и�Z��  �p�"й�"�	 �W�"�Z���R�G_DSBL  ���ˊ���R�IENTTO fZC���A 沽U�`IM_D����O��V�LCT ���Gbԛa�zZd��_PEX�`�7�*�RAT�g d�/%*��UP )���{���������������$PAL򶂷����_POS�_CHU�7����2�>3�L�XL;�p��$�ÿ U�g�y����������� ����	-?Qc@u����Y2C� ��"4FXj |������  //$/6/H/Z/l/~/�Y���.��/�/ςP�/??,?>?P? b?t?�?�?�?�?�?�? �?OO�/�/LO^OpO �O�O�O�O�O�O�O _ _$_6_H_Z_)O;O�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�_����o�m ��� (�"{BPw�m�m ���~�jw8��w ������2�T���p��w���H��t	`����̏ޏ��:��o����� �2���A�  I��j�`� ��������џ�@��@��#�)�Or��1����� 8���, �\Ԡ�� @D7�  ��?���~�q?� ���!D�������%G�  ;�	�l��	 ��xJ젌x����� �<� ���� ��2�H�(��H3k7H�SM5G�22G���GN�3%�`R��oR�d�2�Cf��	a��{�ׄ���������3��¸��4��>���К�����3��A�q½{q��!ª��ֱ� "�(«�=�2������ ��{  �@�Њ���  ���Њ�2��ς�	�'� � ���I� �  y�V���=�������˖ß���  �~y��n @"� �]�<߭˄�����r��N�Д�  '����w�ӰC��C��\C߰��Ϲ��ߤ!^���@�4���/��2�~�B��B�I�;�)�j客z+��������������(� �� -���#�������!��]�9��  q�?��ffaH�Z��� !��������8� ��B��>�|P��}�(� ��P�������\ӯ?��� x� ����<
6b<���;܍�<����<���<�^��*�gv�A)ۙ��脣��F�?fff�?}�?&� ��@��.��J<?�;\��N\��)� ����������� ޤy�N9r]�� �����/&/� J/5/n/�	g/�/�c(G@ G@0~i�G�� G}�� �/??<?'?`?K?�?�o?BLi�B��A �?y?�?|��?K�?ů �/QO�/xO�?�O�O�O<�Om��b��n�t @|�O'_�OK_6_H_�_�3��A��RS�i�Cn_�_j_0O�]?��ooAo,où��Wi���ToC����`CHQo>Jd�x`a�a@Iܚ>�(hA� �A�LffA]��??�$�?���ź�°u�æ�)��	ff��Cϼ#�
�opg\�)��33C�
������<�����nG�B����L�B�s����	0�źH�ۚG���!G��WIY�E���C�+��½I۪I��5�HgMG��3E��RC��j=�~
�pI����G��fIV�=�E<YD �#Zo���
��U� @�y�d���������я �����?�*�c�N� ��r��������̟� �)��9�_�J���n� ����˯���گ�%� �I�4�m�X���|��� ǿ���ֿ���3�� W�B�Tύ�xϱϜ��� ������	�/��S�>� w�bߛ߆߿ߪ߼��߀����=�(�a�L�(�q��)��<��Z������a3�8������a�4Mgu�����a��VwQ�(�4p�+4�]B�B���@p����������UPb	P���QO%x�10[FjR��`�����  C���I4mX��8
O���� ��.//>/d/R/�Rj/|/�/�/�/�/�/�:  2 Fs��gGT�&6��M�eBmp�R�P�aC��3@�_p?�?�?�?�?�?�=�S�OO�)O;OMO�c?��ͫ@@�j��`��`�1�`�^
 TO�O�O�O�O�O_ #_5_G_Y_k_}_�_�_��j�A ����D���$PARA�M_MENU ?�B�� � DEF�PULSE�[	�WAITTMOU�TkRCVo �SHELL_�WRK.$CUR�_STYL`�DlOPTZ1ZoPT�BooibC?oR_DECSN`���l�o �o�o&OJ \n������Q�SSREL_ID�  >�
1��uU�SE_PROG �%�Z%�@��sC�CR` �
1�SS�_HOST !�Z#!X���M�T _����x������L�_�TIMEb �h�~�PGDEBUG�p��[�sGINP_FOLMSK�E�T� \V�G�PGAr� 5���?��CHS�D�TWYPE�\�0� �
�3�.�@�R�{�v� ����ï��Я��� �*�S�N�`�r����� �����޿��+�&� 8�J�s�nπϒϻ�G�WORD ?	�[
 	PR2���MAI�`�3SU�a��TEԀ���	Sd�COLА�C߸�L� �C�~�h�d*�T�RACECTL �1�B��Q }��9 :'���0�ށ�DT Q�B��М�D � � �@U���������������T ��� ����T*��T�T�T�S0���� �����@���f�U 1��@��@�⨐�␅@��@���ԟ��*��Ү�Ҷ�Ң@��R������&�֞�U֦�֮�ֶ�־�����.�����R��	����U����S���������ц�����������Ѫ����������Ѫ��&��.��^�Ѫf��n�О�Ц�Ъ��ж��F�����*��І�Ў������T��G����Ӟ�Ӧ�UӮ�Ӷ��F��N����Ҏ�����i��U�6�>�����>�O��O��O���O��OF�O��O���O��O��O.O
6O>O����3��՞�զ�ծ��
���F��N�'�U�O��O�O&�O.�O*�$O�$O�$O��%�_�Of�On�Ov�OJ~�O��O����^檟�T��T��T��T�F�T��T��T��T���T&$T6T>TP�/�Ԟ�Ԧ�UԮ�Զ��F��N� 9�Ѥ�(O:OLO^O pO�O�O�O�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�P�$Or��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~�f�� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�a��$PGTRACELEN  �a�  ����`��f_UP �����q�'pq p�a_C�FG �uT	s�a p�LtLt�fqwpqz  ��qu4rDEFSP/D �?|�ap���`H_CON?FIG �usW �`�`d�tM��b �a�qP�t؃q��`��`IN~7pTRL �?}�_q8�u�PE�u��w�qLt�q\qv�`LID8s�?}�	v�LLB 1¾�y ��B��pB4Ńqv ��އ؏	�s <o< �a?�� '���A�o�U�w��� ����۟��ӟ��#�	�+�Y�v�񂍯���� ï
��������/�u��GRP 1ƪ���a@�j���hs�aA�
D��� D@� C�ŀ @�٭^��t�q�����q�p�`��.� ���Ⱦ´���ʻB�)�	����?�)�c��a>��>�,��Ϻ��ζ�� =49X=H�9��
����@�+�d� O���s߬�o߼����ߏ  Dz���`
 ��8���H�n�Y��}� �������������4���X�C�|���)���
V7.10be�ta1Xv Aw������!������?!G�>�\=y�#��{3�3A!��@���͵��8wA���@� A�s�@Ls���� ��"4XFXLsApLry��ā��_��@l���@�33q�`�s��k��An�ff�a��ھ���)�x�� �ar�T�n�t�����	t�KNOW_M  |uGvz��SV ��z �r�&����>/@�/G/�a��y�MM�]��{ ���	^u? (l+/�/�',_t@X&Ls����@���%��"4�.N�z�MR
M��|-TU�y�c?�u;eOADBANgFWD~x�STM��1 1�y�4�Garra_]B�2Sem�X�?~s�;Co�2���O�7�3Ante�na_Full @��VODe�qH�� ^OpO�O�O�O�O�O�O !_ __W_6_H_�_l_�~_�_�b�72�<�!4>�_  �<�_�_�N�3�_�_
oo�74 9oKo]ooo�75�o�o�o�o�76�o�o��772DVh�78`�����7MA�0���swwOVL/D  �{�/a��2PARNUM � �;]��u�SC-H*� 8�
����8ω�3�UPD��[��ܵ+�wu_CMP_0r -��0�'�5C��ER_CHKQ�����1�"e�N�`�RqS>0�?G�_MO�?�_��#u_RES+_G�0��{
Ϳ @�3�d�W���{����� ���կ���*�����P��O��8` l�������`��ʿϿ ��`�	���1p)� H�M���phχό����p�������V 1���5�1�!@`y��ŒTHR_IN�R>0/�Z"�5d:�M�ASSG� Z[�M�NF�y�MON_QUEUE ��5X�6Ӑ~  #tNH��U��N�ֲ���ENqD�����EXE�ߌ���BE������O�PTIO������P�ROGRAM %��%��߰���?TASK_I,�>�OCFG ά�x]�����DATAu#��������2� O�?�OTE�U��^�p������:� � ��������������� ~ x ~� �/AS�IN+FOu#� ���Ԕ$ ������
 .@Rdv��� ����/as x�� � ;���ȀK�_�����S&ECNB-�b-&q�&2�/ڝ(G��2�b+ �X,		��=�{���/��@��P4$�0��99)�N'�_EDIT ����W?i?��WERF�L�-ӱ3RGAD�J �F:A�  �5?Ӑ�5Wј6���]!֐��??�  Bz�WӐ<1Ӑ�%�%O�8�;��50!2��7�	�H��l0�,�B=P�0�@�0�M�*�@/�B *�*:�B�O�F�O2��D��A�ЎO�@O	_�,X��%���H�q��O$_r_0_�_���Q@WA��>]�_�_�_o �_o�_�_
o�o.o�o jodovo�o�o�o�o�o �o\XB<N� r����4��0� ��&���J������� ����������x� "�t�^�X�j�䟎��� ʟğ֟P���L�6�0� B���f���������(� ү$������>��� z�t��� Ϫ����� �l��h�R�L�^�DX�	���ώ0�� ���t$ :�L��o�
���ߥ��7PREF S��:�0�0
�5?IORITYX�M6}��1MPDSPV��:
B �UT��C�6�ODUCT���F:��NFOG[@_�TG�0��J:?�HI?BIT_DO�8���TOENT 1��F; (!AF�_INE*������!tcp����!ud��8�!�icm'��N?�X�Y�3�F<��1)�� �A�����0� ����������'  ]D�h�������*>��3���9
BOTf�3?+��F�G/�LC���4�;LFJAB,  ���F!/�/%/7/�5�F�Z@�w/�/�/�/�3&�ENHANCE S�2FBAH+d�?�%;�������Ӓ1��1PORT_N�UM+��0����1_CARTRE�@��q�SKSTyA*��SLGS�������C�U�nothing�?�?OO�۶0TEMP �N�"O�E��0_a_seiban|߅OxߕO�O �O�O�O_�O'__K_ 6_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1U@e� v����������Q�<�u�.IVE�RSI	�L��� �disabl�e'2*KSAVE ��N�	267_0H771|�h���!�/��9�:� !	^�4�ϐ����e��͟ߟ������9�D�C-Å_y� +1���������ő����Ǻ�URG�E� B��r�WF Ϡ��-��9�W�����l:WRUP_DELAY �=�n�WR_HOT �%��7��/p��R_NORMALO��V�_�����SEMI𓿹�����QSKI%Po��97��xf�=� b�a�sυ�H��ʹ��� ���������&��J� \�n�4�Fߤߒ����� �߲���� �F�X�j� 0��|�������� ���0�B�T��x�f����������ãRBT�IF�5���CVT�MOU�7�5����DCRo���� �T�CdE�5E@DA.��@*r�? �>��yH�����č��ğ��H����e����LKUϥ��<
6b<���;܍�>u.��>*��<��AǪP0��� 2DVhz��������,GRDI�O_TYPE  �v��/ED� T_CFG ��-6�BH]�EP)��2��+ ��B�u �/�*��/�? �/%?=�/V?�}?�� �?���?�?�?�?�?O 
O@O*Gl?qO��8O�O �O�O�O�O�O�O�O_ <_^Oc_�O�__�_�_ �_�_�_o�_&oH_Mo l_o�oo�o�o�o�o �o�o�o"DoIho* j������ �.3�E��f� ��� x��������ҏ�*� /�N��b�P���t��� ��Ο��ޟ�:�+���~R'INT 2�R�z�!�1G;� i��{��"���8f�0 ��ӫ����� �M�;�q�W������� ˿���տ�%��I� 7�m��eϣϑ��ϵ� ������!��E�3�i� {�aߟߍ��߱����������A���EFP�OS1 1�!)  x���n# ������������� /��S���w����6� ����l�������= O����6���V �z� 9�] ����Rd� ��#/�G/�k// h/�/</�/`/�/�/? ?�/�/?g?R?�?&? �?J?�?n?�?	O�?-O �?QO�?uO�O"O4OnO �O�O�O�O_�O;_�O 8_q__�_0_�_T_�_ �_�_�_�_7o"o[o�_ oo�o>o�o�oto�o �o!�oEW�o> ���^���� �A��e� ���$��� ��Z�l�����+�Ə O��s��p���D�͟ h�񟌟�'�ԟ� o�Z���.���R�ۯv� د���5�ЯY���}� ��*�<�v�׿¿���� Ϻ�C�޿@�y��e�2 1�q��-�g� ����	��-���Q��� N߇�"߫�F���j��� �ߠ߲���M�8�q�� ��0��T������ ��7���[�����T� ������t�����!�� W��{�:� ^p��A� e �$��Z� ~/�+/���$/ �/p/�/D/�/h/�/�/ �/'?�/K?�/o?
?�? .?@?R?�?�?�?O�? 5O�?YO�?VO�O*O�O NO�OrO�O�O�O�O�O U_@_y__�_8_�_\_ �_�_�_o�_?o�_co �_o"o\o�o�o�o|o �o)�o&_�o� �B�fx�� %��I��m����,� ��Ǐb�돆����3� Ώ���,���x���L� ՟p�������/�ʟS���w�����ϓ�3 1��H�Z������ 6�<�Z���~��{��� O�ؿs����� ϻ�Ϳ ߿�z�eϞ�9���]� �ρ���߷�@���d� �ψ�#�5�G߁����� ��*���N���K�� ��C���g����� ����J�5�n�	���-� ��Q���������4 ��X��Q�� �q���T �x�7�[m �//>/�b/� �/!/�/�/W/�/{/? �/(?�/�/�/!?�?m? �?A?�?e?�?�?�?$O �?HO�?lOO�O+O=O OO�O�O�O_�O2_�O V_�OS_�_'_�_K_�_ o_�_�_�_�_�_Ro=o voo�o5o�oYo�o�o �o�o<�o`�o Y���y�� &��#�\��������?�ȏ����4 1� ˯u�����?�*�c�i� ��"���F����|�� ��)�ğM�����F� ����˯f�﯊���� �I��m����,��� P�b�t������3�ο W��{��xϱ�L��� p��ϔ�߸������ w�bߛ�6߿�Z���~� ����=���a��߅�  �2�D�~�������� '���K���H������ @���d����������� G2k�*�N ����1�U �N���n ��/�/Q/�u/ /�/4/�/X/j/|/�/ ??;?�/_?�/�?? �?�?T?�?x?O�?%O �?�?�?OOjO�O>O �ObO�O�O�O!_�OE_ �Oi__�_(_:_L_�_ �_�_o�_/o�_So�_ Po�o$o�oHo�olo�o<ۏ�5 1����o �o�olW��o�O �s���2��V� �z��'�9�s�ԏ�� �������@�ۏ=�v� ���5���Y��}��� ��۟<�'�`������ ��C���ޯy����&� ��J����	�C����� ȿc�쿇�ϫ��F� �j�ώ�)ϲ�M�_� qϫ����0���T��� x��u߮�I���m��� ���������t�_� ��3��W���{���� ��:���^�����/� A�{����� ��$�� H��E~�=� a�����D/ h�'�K�� �
/�./�R/�� /K/�/�/�/k/�/�/ ?�/?N?�/r??�? 1?�?U?g?y?�?O�? 8O�?\O�?�OO}O�O QO�OuO�O�O"_t6 1�%�O�O_ �_�_�_�O�_|_o�_ o;o�__o�_�oo�o BoTofo�o�o%�o I�omj�>� b������� i�T���(���L�Տp� ҏ���/�ʏS��w� �$�6�p�џ������ ���=�؟:�s���� 2���V�߯z�����د 9�$�]��������@� ��ۿv�����#Ͼ�G� ����@ϡό���`� �τ�ߨ�
�C���g� ߋ�&߯�J�\�nߨ� 	���-���Q���u�� r��F���j����� �������q�\���0� ��T���x�����7 ��[��,>x ����!�E� B{�:�^� ����A/,/e/ / �/$/�/H/�/�/~/?��/+?�/O?5_GT7 1�R_�/?H?�?�? �?�/O�?2O�?/OhO O�O'O�OKO�OoO�O �O�O.__R_�Ov__ �_5_�_�_k_�_�_o �_<o�_�_�_5o�o�o �oUo�oyo�o�o8 �o\�o��?Q c���"��F�� j��g���;�ď_�� �������ˏ�f�Q� ��%���I�ҟm�ϟ� ��,�ǟP��t��!� 3�m�ί��򯍯��� :�կ7�p����/��� S�ܿw�����տ6�!� Z���~�Ϣ�=ϟ��� s��ϗ� ߻�D����� �=ߞ߉���]��߁� 
���@���d��߈� #��G�Y�k����� *���N���r��o��� C���g��������� ��nY�-�Q �u��4�X��|b?t48 1� ?);u��/ ;/�_/�\/�/0/�/ T/�/x/?�/�/�/�/ [?F???�?>?�?b? �?�?�?!O�?EO�?iO OO(ObO�O�O�O�O _�O/_�O,_e_ _�_ $_�_H_�_l_~_�_�_ +ooOo�_soo�o2o �o�oho�o�o�o9 �o�o�o2�~�R �v���5��Y� �}����<�N�`��� ������C�ޏg�� d���8���\�埀�	� ����ȟ�c�N���"� ��F�ϯj�̯���)� įM��q���0�j� ˿��ￊ�Ϯ�7�ҿ 4�m�ϑ�,ϵ�P��� tφϘ���3��W��� {�ߟ�:ߜ���p��� ����A����� �:� ����Z���~���� �=���a���� ������MASK 1���������?XNO  ����~ MOTE  �  N_CFG� �Y����P?L_RANGUP�����OWER ���� �A���*SYSTEM�*P�V9.304�4 �1/9/2�020 A ��g ���REST�ART_T  � , $FLA�G� $DSB_�SIGNAL� �$UP_CND�4P��RS232�r � $�COMMENT �$DEVI�CEUSE4PE�EC$PARIT�Y4OPBITS�4FLOWCON�TRO3TIME�OUe6CU�M�4AUXT��5INTERFACs/TATU�X�SCH t $OLD_y�C_SW 'F�REEFROMS�IZ �ARGE�T_DIR �	$UPDT_M�AP"� TSK_wENB"EXP:*z#!jFAUL �EV!�RV_D�ATA�  �$n E�   �	$VALU�!� 	j&GRP_ �  {!A�  2 �S�CR	� ��$ITP_�" �$NUM� OU�P� �#TOT_A�X��#DSP�&J�OGLI�FIN�E_PCd�ONmD�%$UM�=K5 _MIR1!4�PP TN?8APL"G0_EXb0<$�!�� 814�!PGw6BgRKH�;&NC� �IS �  �2T�YP� �2�"P+ Dxs�#;0BSOC�&�R N�5DUMMY�164�"SV_C�ODE_OP�S�FSPD_OVR5D�2^LDB3�ORGTP; LEbFF�0<G� OV5;SFTJRUNWC!�SFpF5%3UFR�A�JTO�LCH�DLY7RECO1VD'� WS* �0��E0RO��10_~p@   @��}S NVERT"�OFS�@C� "F�WD8A�D4A�1EN�ABZ6�0TR3�$1_`1FDO[6MOB_CM�!FPB� BL_M��!2hRnQ2xCV�"' } �#2PBGiW|8AMz3\P0��U�B�__M�P��M� �1�AT$CA�� �PD�2�PHB�K+!:&aIO�4 �eIDX+bPPAj?a$iOd7e�U7a��CDVC_DBG "�a;!&�`�B5�e�1�j�S�e3�f�@ATIO� ���AaU�c� �S�AB
0Y.#0�D��X!�� _�:&SUBC�PU%0SIN_RS�T, 1N|�S�T�!�1$HW_C�1�"]q.`�v�Q$�AT! � �$UN�IT�4�p�pAT�TRI= �r0CY{CL3NECA�b�L3FLTR_2_�FI9a7�c,!L�P;CHK_�S�CT>3F_�wF_�|8��zFS+�R�rCHAGp�y��R�x�RSD�@'�1E#�&7`_T�XPRO��`@S�EMPER�_0�3Tf�]p� xf��P�DIAG;%?RAILAC�c4r�M� LO�0�A�65&�"PS�"�2 -`�e��SPR�`S.  ��W�Ctaf	�CF�UNC�2�RINS_T.!(�w�L�� S_� �0�Pp�� 	d��WARL0~bCBLCUR���єAʛ�q͘ƘDA`�0���ѓʕLD  @,a3��!��8�3��TID�S��!� $?CE_RIA !5+AFDpPC~��@��T2 �C9#�b{Q�OI�pCVDF_LaE��#0(!�LM�S�FA�@HRDYO,L1	PRG8�H��>1�(�ҥMULSE� =#Sw3��$J�JJ6BKGFKFAN?_ALMLV3R��WRNY�HARDH�0+&_P "��2Q�Ȏ�!�5_�@:&AU��Rk��TO_SBRvb��� ƺ�pvc|�޳MPINF�@��q�)���REG�'d~0V) 0R�C�1DgAL_ \2FL�u�2$MԐ(�#S�d�P� `�g�CMt`3NF�qsONIP�qpEIPP �9a$Y��! ��"�!� ��o3EGP��#@��AR� �c�52������|5AXE�'ROBn�*RED�&WR�@2�1_=��3SY�0�t�0_�Si�WRI�@�ƅpST�#��0*@� �q	���3��� �B� �A��3�D�PO�TO�� �@AR�Y�#��!��d�!1F�I�0�$LIN]K��GTH�B ST_���A��6�"N/�XYZ+"9�7G�'OFF�@�.�"�%��B� l����A3$ ��FI�p���h4�4l��$_Jd��"(B�,a������8@�"q������C�k6DUR��94�TURT�XZ�N����1Xx��P��FL/�@`s��l�P��30�"^Q 1� K
0	M:$�53]q7�SuD�Sw#ORQɆ�!��P���Q7��0O[�ND��=#�!#�1OVE8��M���R�� R��Q!P.!P! OAN}q	�R���� 990� �brJ9V`����v�!ER1
��	8�E�@n D�	A��p�嘕Ă���v�AX�C�"� �`�q�s�� �0~3�~F�~e�~�~E�~1��~Ҡ {Ҡ�Ҡ�Ҡ�Ҡ �Ҡ�Ҡ�Ҡ�Ҡx�!)DEBU}s$x���삼!R*�CAB�a8A2V`|r 
�"�c���% �Q7�7�173�7 F�7e�7�7E�p������LAB��q��yp�cGRO�p4��}��PB_ҁ  ��̓��ð�6�1���5���6AND��8p �a3���-G �Q�����AH�PH�p2�NT8d��Cs@VEL؁��}A��F�SERV9Es@�� $����mA!�!�@POR }�KP�иA���@����	��$�BTREQ�
�CH��@
�GƄ�2	�Eb��_ � lb��Q�ERR��RI�P�@�NFQTOQ�� L�P}��YVĀG�E%��\���BRE� G ,�A�EP
��RA�Q 2 �d�R7c�U�@ ��$F ׂ��m�UOC��P � 8[COUNT����A�SFZN_wCFG�A 4�p%��rT\zs�a�#`p�Jp�q��&c�� �� MGp+���`�`�OGp�eFAq����cX8еk�ioQH��'ѴDp8�Pz�?��SHELA�-b� 5��B�_BAS\RSR$�`�2�S��L�!p�1�W!p2Dz3Dz4�Dz5Dz6Dz7Dz8�WqROO���P�f1�NL�� �AB�C�
�"pACK�&IN�PT+�W�U��	�k���y_PU8�~�|�OU�CP��%�s�Vl����YTPFWD_�KARKQ-�:PREĿD�P����QUE$�Ā9 )���~���IU��#s/���@�/�SEM1ǆ1��A�aSTY�tSO����DI�q��Qc���X��_TM9�MA�NRQ �/�END���$KEYSWITCH2�G�����HE)�BEATM6z�PE��LEJR����0x�UF�F��G�S~�DO_HOM���Oz��pEFPR���SbJі��uC��Ox��7P�QOV_M��<}�c�IOCM����1��tHK��# D,�&�a`U2R���M��a�r +�FOR�C*�WAR��O}M��  @�$T�㰰U��P�1��g���3��4�1�B�P�OW�Lz��R%�U�NLO�0T�E�D��  �SNuP��S.b 0N��ADDa`z�$S{IZ*�$VA�0~�UMULTIP�r����Az� � $��ƒ����SQc�1CFPv�F'RIFr�PSw����ʔf�NF#�ODBUx�R@w������F��:�IAh�����������S"p�� �  �cRTE���SGL.�T�x�&�C`Gõ3a�/�STM�T��`�P����BW<9 0�SHOWh�q7BANt�TPo���@E������@V�_Gsb �$PaC�0�PoFBv�-P��SP��A�p����`VD��rbw� �+QA002D .ҝ�6ק�6ױ�6׻��6�54�64�74�8*4�94�A4�B4و� 6ׇ17�}�6�F4�  ��@�����Z����t�U1��1��1��1��U1��1��1��1��U1��1��23�2@�U2M�2Z�2g�2t�U2��2��2��2��U2��2��2��2��2��2��33�����M�3Z�3g�3t�3���3��3��3��3���3��3��3��3���3��43�4@�4�M�4Z�4g�4t�4���4��4��4��4���4��4��4��4���4��53�5@�5�M�5Z�5g�5t�5���5��5��5��5���5��5��5��5���5��63�6@�6�M�6Z�6g�6t�6���6��6��6��6���6��6��6��6���6��73�7@�7�M�7Z�7g�7t�7���7��7��7��7���7��7��7��7���7���VPv�U�B �@�09r�
�����A x e�0R���  �B�M�@RP�`�4Q_��PR�@[U�AR��DS�MC��E2F_U8��=A��YSL�P�@ �  �ֲ>g��������iD��VALU>e�pL�A�H=FZAID_L���E�HI�JIh�$FI�LE_ ��D�d$�ǓB�XCSA�Q� h�0!PE_BL�CKz�.RI�7XD_CPUGY!�GY�Ic��O
T�PY.��R � � PW�`�p���QLAn��S�Q�S�Q�TRUN_FLG�U�T�Q�T@J��U�Q�T�Q�UH�p�T`�T��T2L��_LIz�  ]�pG_OT��P_EDIU�X /`�`7c ?bة�p�BQh�����TBC=2 �! �%�>�0�P��a�7aFTτ�d.݃TDC�PA�N`��`M�0�f�a�gTHD��U��d�3�gR�q<�9�ERVEЃt�݃t	��a�p�` "X -$EqLENЃRt݃Ep�pcRAv��Y@W_A�tS1Eq�D2�wMO$?Q�S���pI�.B`�A�y�4Ep�{DE�u���LACE �CCqC�.B��_MA�p�v��w�TCV�:��wT,�;�Z�P�Ҡ�s��~��s��J�A��M����J���u)ā�uQq2ѐ����݁�s�JK��V�K������	���J�����JJ�JJ�AAL�<��<��6��:�5�cm�N1�a�m�,��DL�p_�\�Ű�ApCF
�#{ `�0GROU�@(J�Բ��N�`C^�Ȑ?REQUIRrÀ�EBUu�Aq��$T�p2"��Bp薋a�	��d$ \?@qhA�PPR��CLB
u$H`N;�CLO}`"K�S�e`��u
�aI�% �3�M�`�l���_MG񱥠C� �"P����&���BR=K��NOLD����RTMO6a�ޭ��	J6`�P>��p��p@��pZ��pc��p6+��7+�<�B����e&G� �lr����<����PATH����@����qx�����%0A��SCAub��<���INDrUC�p�q�-C�UM�Y�psP����A q/ʤ�/��E�/�PAYLOA��J2L�0R_A	N�ap�L�Pz�v�j������R_F2LS3HRt��LO{�R�������ACRL�_�q�����b�d�H��@B$H��"�FWLEX>���J�f' P(��o�o+�p�>�Du( :Qcv�p����fe�0�po��|F1��� -������]�E��*�<�N�`�r� ����4�Q�������A�@c���ɏۏ���T��2�X:A;����� ����)�;�?�H�@6�Z�c�u�����P=���) ��`��˟ݟ��`�0ATF�𑢀E�L��(a��J�(v��JE۠CTR���A�TN�1�HA_ND_VBB>�ܯ@�* $��F24���d�CSWR�����+� $$M �����0ˡ�ڡ������A�@g����AD)��A���@˪A٫AA� ��`P˪D٫�D�PȰG�P�)S�Tͧ�!ک�!N�DY�P9����#%��Fp ���Ѫ���i����������P3�<�E�N�W��`�i�r�RD���,c ��ԓ� n�x�5m��1ASYMص.@�ض+A������_`��	���D@�&�8�J�\�n�Ju��&��ʧC�I��S�_V�Io�Hm��@V_�UNVb�@
S+��J �"RP5"R��&T��3T WV�͢���&��ߪU���/�7�<ѓ`HR`ta-��QQ�1�DI��O�T���PN��. ; *"IAA*���$aG�2C2cJ���`]`I��P / �� �ME��� Mb�R4AT�PPT@�@� ��ua���PАl@zh�a�iT�@��� $DUMMY}1E�$PS_D�RFॐ$�fn3�FLA��YP����b}c$GLB_T��Uuu`1�����EQa0 X(����ST����SBR��PM21_V��T�$SV_ER��O�_@KscsCLpKrA���O'b�PGL�@E�W��1 4��a+$Y|Z|W�s�D���AN`vU�u�2 ��N�p�@w$GIU}$�q 1_�s�p���3 L���v^B}$�F^BE�vNEARʖ�NK�F8���TA�NCK�����JsOG��� 4��$JOINT��x� ��qMSET��5  �wE�H�� �S��Q�� ��6��  MU��?����LOCK_FOx����PBGLVH�GL�TEST_sXM>���EMPt�����r̀$U�Гr��22���s,��3���Ҁ,�1MqC�E���sM� $KA�R��M�STPDRqA�pj�a�VEC�Ь{�e�IU,�41�H=EԀTOOL㠓�V�RE��IS3����6N�A�ACH���5��O�}c�d�3���pSI.� � @$RAIL__BOXE��ppoROBO��?�pq?HOWWAR*��<�`�ROLM�bB����S��
�5���O�_F� !ppHT'ML5�Q������2�pڑ��7m�+�R��O��8���v�z���sOU��9 tpp(�14A��̀��PO֡%PIP��N��
�ڑ�S�,�����CORD�EDҀް̠5�XT���q)�S� O4` �: D pOBP!"Ҁ{�j��cp�j�^@$SYSj�A�DR#�Pu`TCH�� ; ,��E�N�RZ�Aف_�t�״�>��PVWV�APa< � �p��r�UPREV_�RT]1$EDI}T�VSHWR��7v;���q�@D�_`#R�+$H�EADoA�Pl�A�$�KE�q�`CPS�PD��JMP��Ld�U=�R��d=r�TO�϶I�S#Ci�NE��$_TIC)K�AMX��q��{HN-q> @t�8�����_GP���[�STYѲ�LO�q�s��Ҩ�?�
��Gݵ%$���t=:7pS !$Q��da�e!`�fP�0�S�QUd� ��b�ATE�RCy`|�S�@ �pCp�����d�%Oz`mcO�I�Z�d�q�e�aPR`M��a8����PUQ�H�_DO=�ְXS:��K�VAXIg�f�1�UR� ��$#��Е��� _����EET��Pۂ���5f��F�7g�A�!�1��d9�2;]�T{SR|Al�� ����#��5��#� �#�)#�)i�>'i� N'i�^&{����){���$�2��C����C��WOpiO{O�DIaSSCp� B hppDS�(�k��`SP`�A	TL �I���¼b�ADDRES��B�'�SHIF��"�_W2CH#��I&p���TU&pI� �C��CUSTOT��qV��IbDȲ,��0
�ߠqV�X�R`E \������f�7��tC��#	���F��irt�TXSCREEl��F�P��TINA�s�p��t�����0G T��fp,⧱ eqBp&uᦲu�$#�RRO'0R���}�!����UE��H ���0���`S�q��RS	M�k�UV����V~!�PS_�s�&C�!�)��'C��Cǂz"� �2G~�UE�4Ipbvr�&8�GMTjP�LDQ��Rp���B�BL_�W�`R`JS �C>2O�qJ2�LE�U3"�T4RwIGH^3BRDxt��CKGR�`�5T�W��7�1WIDTH��H������a��7�UIu�EY��QaK d�p��A�J�
�=4�BACKH��b4�5|qX`FOD�G�LABS�?(X`I<�˂$UR(�9@����0^`H4! L 8�QR�_k��\B_`R�p͂�����HB)O�R`M��w0�Uj0�CRۂM�LUqM�C��� ERV���p�0P<��4NV`��GE=B#���]�t��LP�E��E��Z)�Wj'Xz'XԐ&Y5*$[6$[7$[8	R��@�3�<���fԑŁ�S��M�1USR��tO <��^`U��r�rFO
�rP�RI��m����PT�RIP�m�U�NDO��P�p ��`m�4���#����� QWB�P7�G �s�Tf�H�RbO	S�agfR��:">c��.qR��s�~�b*�� #�UQ.qS�o�o�#8R)�>cOFF���p�T� �cOp �1R�t/tS�GU��P.q��JsETwn�1SUB*� f�_E_EXE��V��v>cWO>� U�`^g��WA'��P�q�!@� V_DB��s�p��PT�`
�V0�Q�r��OR��u'RAU��tT�ͷr�q_���W |%��͸OWNA`޴$GSRCE � ��D��<\��MPFIA�p��ESPD����� �C���Gƒ] +�5��!GX `�`�r޴�n��COP�a$��C`_w������rCT�3�q���qƒ����@� Y"SHADOW�ઓ@�?_UNSCA��@���4M�DGDߑ��E�GAC�,��PG��Z (0NOX�@�D<�PE�B��VW� �G���![o � ��VEE#��ڒANG�$��c�薴cڒLIM_X �c��c� ����#`��`� 퐾�VF� ��s�VCCjв�\ՒC{�RAlצ���\RpNFA��Z%�E��Z`G� f^0[�C`DEĒ��� STEQ1���@ �ꁻ@I��`+0���p�`����P_A6��r���K��!]�# 1Ҡ�����\�ȫсCPC�@]�DRIܐ\�͑V#Ѐ����D�TMY_UBY�T���c��F!���bY��$���P_V��y��LN�BMQ1�$��DEY��EXX�e��MU��X�M� US�!���P_AR����P� ߖG��PACIr�ʐf�ᔀ���c�´c���#�EqB��a.2B���Ч^ ܀GΐP����� C�R~``�_ �0�@3!�1zr	�e�R�SW��p�00��$S�6�O�Q�1A� XӚ#�E�UE��00�)�D�HKJ�`�@�p���U� �EA�N�ٖp�pXՆ`C�MwRCV�!a ��@UO��M�pC�	��8s����REF*7
� �������/��P��@�@��@��b��֗�_Y� �ژ��ۣ��Q$3������C��$b �����%���Q��$GROU� �c���d��ʠ]��I2^00��U` 0_�IX,�o � ULա`���C&�rAaB�?�NT����$����A���Q��K�L����õ��A����Q��T a$c �t�`MD�p8�HUح��SA��CM�PE F  _��Rr�p@����X<S	�VGF/�b#_d, &�@M�P^0۰UF_C !���z �ROh0"+��p�@���0C�UREB����RI��
IN �p�����d��d�,�ca�INE�H�y��0V�a-�걗�3�W�������C��i�LO�}�z�@0�!�QNSI��݁����c$&�c$&.�X_PuE-YW+Z_M�ڒW�I�$�" �+�R�'rRSLre� �/�M
`�RE�C7�Gd�۰�� �ҭ�q����u��� �������S_P�V�nP  �VIA�vf �~pHDR��p7pJO�P��$Z_UP�=�a_LOW�5�1tJ�dA��LINubEP?�tc_i�1�1����@�G1@��V�xg� 5X�PAT�HS� X�CACH $�]E��yI�A��*{�C)�ID3FA�EsTD�H��$HO�p"O�b@�{�d6�F������p�PAGE��䁀VP�°�(R_'SIZ��2TZ3�-X0�0U�q�MPRZ���IMG���AD�Y�MRE��R7W�GP��8�p��AS�YNBUF�VR�TD�U�T7Q�LE�_2D-��U��`C�ҡU1��Qu��UEwCCU��VEM��x]EDb�GVIRC�Q`�U�S�B�Q�LA�þp�NFOUN_�D�IAG�YRE�XYZ�cE�WѴh8ȳdpqa`T��2�IM��a�V|be��EGRA�BB��Y�a�LE%Rj�C4���FC-A��6504x��7u$��pBE��h��`�CKLAS_@l�BA��NN@i  G��T��S�@ݲմ$BAƠwj �!q�eb��u�TYSp�H����2��I��t:b�f��B)�EVE����PK���fx6��GI�pNO��2��ER�rHO����k � ���
8��Pi�S�0ޗ��RO>��ACCEL?0=�-��VR_�U7@�`���2�p��AR��P�A��̎K�D��RE�M_But �1S'_JMX �l�t�$SSC�Uk��p#���QN@m � ��S�P�NS���L�EX�vn T�E�NAB 2�W@��F7LDRߨFI�P��t�ߨ(Ğ��"P2>HFo� ���V
Q MV_PI ��8T@󐉰�	F@�Z�+�#��`8�8#��GAB�Ε�LOO��JCqBx��w"SCON(P�PLANۀ�Dp��3F�d�v�9PէM ��Q ;����SM0E� ɥ�8ɥWb72$`d<�8T��,`RKh"^ǁVANC�� �0�R_Ou N@p ( �-#<#c��c2?B�R_A/�N@q 4 ������`	�^����r hn���1^�&'OFF`|�p�`��,�`�DEA�
�P,`�SK�DMP6VIE��2q w��@��>�rs < {���D�4���r{7��D�����u�CUSTz�U��t $G��TIT1$P9R\��OPTap �O�VSF�йsu�p��0`r&���SMEOwvI�|�ĄJ������eQ_WB��w�I���� @O3�@�7XVRxxmr���T��$�ZAB=C��y op��t��)�
���ZD$��CSCH��z L u����`�2�%PC ��7PGN ��<��A��_FUNH��@o7ZIPw{I��KLV,SL��~��_ZMPCF��|���E����X�DMY_LNH�=�D�� ��?} $�A� ^]�CMCM� C,S�C&!��P�� O$J���DQ��������������_0�Q,2����UX�a\�UXEUL��a�� ����(�:�(�J���FTFL��w����~�0+�6�Џ��Y@Dp  _8 $R�PU���> EIGH����?(�iֱ�@@��et�� �a�����$�B�0�0@�	�_SgHIFD3-�RVV`�Fcв�	$5��C �0��&!������b�
�sx�uD�TR���V̱��SP9H���!� ,�������� �4A�RY�P��%���~��%��@!�%!���H�(UN0���"�@2�����s��q0GSPDak����P��O��`��0�ĳ��}"!NGVER`q7 iw+�I_AIRPUR�GE  i C i/�F`E�Tb�� �+1h2ISO�LC  �,�"� � �!�%��P+Y�_/*OB��Dm��?@�!H771  34 n?�?�9� `�E/#�)�x� S232�� �1i� L�TEk@ PEN�DA�341 1D�3<*? �Maintena�nce Cons� B�? F"O,D?No UseMJO OnO�O�O�O�O2�2GNPO;/" 19%��1CH=� ��.P		9Q_!�UD1:___RSMAVAIL/��/%�A!SR  �+��H�_�P1�oTVAL.&����P(.�YVL�}� 2�i�� D?�P��/`oVPNo�o rci�o�g�o�o�o�o �o*,>tb �������� �:�(�^�L���p��� ����܏ʏ ��$�� H�6�X�~�l�����Ɵ ���؟�����D�2� h�V���z�������� ԯ
���.��R�@�b� d�v�����п����⿀��(�N�<�r�i��$SAF_DO_PULS. j>ap�����CA� �/%��&0SCR ��`X���`�`
	14�1IAIE���b vo$�6�H�Z� l�~�ߢߴ������߬���HS��2�%�����d1�(�8�8rb��� @�"k� }���T�h� J`���_ @��T7 �����#�0�T D��0�Y�k� }��������������� 1CUgy�O<�Ef������  �5;�#o�� 1p�U��
�t��Di��������
  � ��*������gy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7O<A���`OrO�O�O�O�O �O�O�O?O�_._@_ R_d_v_�_�_�_�_�Q _�R0MJTo !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ JO��'�9�K�]�o� ������_ɟ۟��� �#�5�G�Y��_�U�_ �ҙ�����ϯ��� �)�;�M�_�m����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B�T�f�;�?�q߮� ����������,�>� P�b�t�������������������Y��	123456781�h!B!�)���F����� ������������  ��;M_q�� �����% 7I[l*��� ����//1/C/ U/g/y/�/�/�/n� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? O�/)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_O_�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�op_ �o�o�o/AS ew������ ���o+�=�O�a�s� ��������͏ߏ�� �'�9�K�]������ ����ɟ۟����#� 5�G�Y�k�}�������"��s�կ�w����0�L�CH  �Bpw�   ��=�2�� }� =�
���  	�o�ί���ǿٿ���r���� ��@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖ�%Ϻ��� ������&�8�J�\� n����������� ���"�Q�*������;�<M���D���  �]�w�*��Z򛱛�t  �d�����*�`*��$�SCR_GRP �1*P�3 � �*�� 6�	 �� 
��<�+*�'pUC|@��y�yD� W�!��y�	M-10�iA/7L 12�34567890ڙ�� 8��M1T� � �
�	L���	Č� N 
���Y���y�
M_	P������ ,��#H�
 ���1/�@A/g/y/H�ߙ! T/�/P/�/3��+���/B�S��,?*2C4r&Ad�R?  @0j5N?�7?��7&2R���?}:&F@ F�`�2�?�/�?�?O O-OSO>OwObO�O=�j1�2�O�O�O�O�DB��O�O;_&___J_�_ n_�_�_�_�_�_o�_ %o�5j�eSgxo6����uo�o�b�1�B̃|3�oh0�4j9j9B� w�$Y̯@HtA�Nhcu�/�%Ipp�drsq ����z�q�x� �.� (&�*�2� D�V�oz�e��������ECLVL  Ψ���iqpQ@���L_DEFAU�LT �����փHOT�STR�qq��MIPOWERF���H���WFDO�� �RVENT 1ɁɁ�� L!DUM�_EIP�����j�!AF_INEx‧���!FT}��֞����!-/� ���F�!RP?C_MAING�)�q�5���Y�VISb��t����ޯ!TP&ѠPUկ��dͯ*��!
PMON_POROXY+���e��v��D���fe�¿!�RDM_SRV�ÿ��g���!R�,*ϑ�h��Z�!
�[�M����iIϦ�!RLSYNC�����8����!R3OS|���4��>��!
CE�MTC�OM?ߓ�k-ߊ�!=	S�CONS�ߒ��ly���!S�WA'SRCݿ��m��"�;!S�USB#�n�n�!STMC��o]����� ѳ����,���P�V��ICE_KL ?�%d� (%S?VCPRG1S�����2�������o����4������5��6;@��7ch��H���9���� %��������0 ����X�����- ���U���}��� � /���H/���p/ ���/��F�/��n �/��?��8?�� �`?��/�?��6/�? ��^/�?��/X�j�� q���#OhO��lO�O{O �O�O�O�O�O�O _2_ _V_A_z_e_�_�_�_ �_�_�_�_oo@o+o doOo�o�o�o�o�o�o �o�o*<`K �o������ �&��J�5�n�Y����}���ȏ���^�_D�EV d���MC:�4����GRP 2�d���bx 	�� 
 ,V� ȡ�s�Z������� �����ߟ��@�'� 9�v�]�������Я��P��۫Y���� ܯI�1�4�]���j��� ��˿F�Ŀ��%�7� �[�B��f�xϵ�� !���A����ۿD�+� h�Oߌ�s߅��ߩ��� ��
���@�'�d�v��	y��^������ ����%��I�0�Y�� f�����8���������@��3��T7]�e �����)��
 �.@�dK�o@��!�9�� �!/G/���R/�/�/ �/�/�/"�/�/?? C?*?<?y?`?�?��? �?�?�?�?�?-OOQO 8OaO�OnO�O�O�O�O �O_�O)_;_"___�? �_�_L_�_�_�_�_�_ o�_7oo0omoTo�o xo�o�o�o�o�o! x_E�oU{b�� ������/�� S�:�w�^�p�����я��d �X�ZI�6 r��@�Z��0�+A�����dBj?BA�=��������B����AZ.�AĊ��+�A.�Q��B����5\���i6�A�u���'����%�Ꮛ�%PE�GA_BARRA�_ESTEIRA|����X�T����?=��=X���7
�?�>��A����������&���������Ax�P��f��U��'A�j������B�:��<�3����jB]+����T��%�T���d��ʐ���>�pc?���7�ԳT@�6��A�_���0n�����·�Ak���۸I�K9FA��G����B�!v,�-��C�3�����pBM�>�#�b�(�Y��������HX�?�L!���Q�B����AJ���Xk�@fD3���O�A��������Yw����.B�B��;��CH��z�B�?@���6���-Ϙ������n��=]����V@��?,������� վ��e�Ak�������OY�A������AB�J��;%�C$4�aƿBXZ9濠��
���ߘ�Ţ��� �ԭ(��^_���-\¯ԡ���گ���+����@��������ߔ�ᢧۙ�*נ�6��>�ԯb���zװ>
��BM��sﰲ�x�U<�߯�7@6|=���P�$�6��� N�@���b�G���L�}��������x7��~�K@���V��+A>r�r�F���������Y@+�@�<B���|�A�F�����B)���,o�?ɇ��~0��0~6��Z� Q�杚��������A�ߍ�]ܖA�?���������2[����>��ȥA��=�����NB ��$�w?�dj��to�7\�
`�.�%��Z�����A������*�@Ve�B� ������YN�#�B�D�	���9A����gB#
q�3���C4#��,??[BVM����COLOCA?_PRENS�����&//J/8/n/ \/~/�/�/�/�/ �/ ??D?2?T?�/�/ �?�/z?�?�?�?�?O 
O@O�?gO�?0O�O,O �O�O�O�O�O_ZO?_ ~O_r_`_�_�_�_�_ �_�_2_oV_�_Jo8o no\o�o�o�o�o
o�o .o�o"F4jX ��o��~�z� ��B�0�f����� V�����Џҏ��� >���e���.������� ��̟Ο���X�=�|� �p�^���������ȯ �D��T��H�6�l� Z���~�����ۿ��� Ϡ��D�2�h�Vό� ο���|�����
��� �@�.�dߦϋ���T� �߬���������<� ~�c��,����� �����D�)�;���� ��\������������ @���4"DFX �|����� �0@BT�� ��z��/�,/ /</���/�b/�/ �/�/�/?�/(?j/O? �/?�??�?�?�?�? �? OB?'Of?�?ZOHO ~OlO�O�O�O�OO�O >O�O2_ _V_D_z_h_ �_�_�O�__�_
o�_ .ooRo@ovo�_�o�o fo�obo�o�o* N�ou�o>��� ����&�hM�� ���n���������ȏ ��@�%�d��X�F�|� j��������,���<� ֟0��T�B�x�f��� ޟï��������,� �P�>�t�����گd� ο�����(��L� ��sϲ�<Ϧϔ��ϸ� ������$�f�Kߊ�� ~�lߢߐ��ߴ���,� �#�������D�z�h� ��������(��� 
�,�.�@�v�d����� �� �������( *<r�����b� ���$z� q�J����� �/R7/v /j/� z/�/�/�/�/�/*/? N/�/B?0?f?T?v?�? �?�??�?&?�?OO >O,ObOPOrO�O�?�O �?�O�O�O__:_(_ ^_�O�_�_N_p_J_�_ �_�_o o6ox_]o�_ &o�o~o�o�o�o�o�o Po5to�ohV� z����(�L �@�.�d�R���v��� ���$�����<� *�`�N���Ə���t� ޟp����8�&�\� ����L�����گȯ ����4�v�[���$� ��|�����ֿĿ�� N�3�r���f�Tϊ�x� �Ϝ����������� ��,�b�P߆�tߪ��� ��ߚ������(� ^�L���ߩ���r��� �� �����$�Z��� ����J����������� ��b���Y��2� z�����: ^�R�b�v� ���6�*// N/</^/�/r/�/��/ /�/?�/&??J?8? Z?�?�/�?�/p?�?�? �?�?"OOFO�?mOO 6OXO2O�O�O�O�O�O _`OE_�O_x_f_�_ �_�_�_�_�_8_o\_ �_Po>otobo�o�o�o �oo�o4o�o(L :p^��o�o� � ��$��H�6�l� ����\�ƏX�֏�� � ��D���k���4� ������ҟ���� ^�C����v�d����� ����ί��6��Z�� N�<�r�`��������� �󿪿̿���J�8� n�\ϒ�Կ�������� �������F�4�j߬� ����Z��߲������� ���B��i��2�� �����������J�p� A����t�b������� ����"�F���:�� Jp^������ � 6$Fl Z������� /�2/ /B/h/��/ �X/�/�/�/�/
?�/ .?p/U?g??@??�? �?�?�?�?OH?-Ol? �?`ONOpOrO�O�O�O �O O_DO�O8_&_\_ J_l_n_�_�_�O�__ �_o�_4o"oXoFoho �_�_�o�_�o�o�o �o0T�o{�oD �@�����,� nS�����t����� ����Ώ�F�+�j�� ^�L���p�������ܟ ��B�̟6�$�Z�H� ~�l����ɯۯ���� ����2� �V�D�z���������$SE�RV_MAIL + �����ʴ�OUTPUTո��@ʴRoV 2j�  㰧 (r����x��=�ʴSAVE����TOP10 2�� d 6 rƱ���϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t������n�YPY��FZN_CFG f��=��J���?GRP 2��g�� ,B   A� =�D;� B� �  B4=��RB21I�HELL��f�e�)��*�=�����%RSR����� �&J5G� k������.?�  ��/�>/P/"\/ ��X/z"{ �U'&"2��dh,g-�"EHKw 1S �/ �/�/�/#?L?G?Y?k? �?�?�?�?�?�?�?�?�$OO1OCO?OMM� S�ODFT?OV_ENBմ��e��"OW_REG�_UI�O�IMI_OFWDL~@�N��BWAIT�B �)��V��F�YwTIM�E��G_�VA԰_�A_UNcIT�C~Ve�LC�@WTRY�Ge�ʰ�MON_ALIA�S ?e�I%�he��oo&o8oFj�_ io{o�o�oJo�o�o�o �o�o/ASew "������� �+�=��N�s����� ��T�͏ߏ����� 9�K�]�o���,����� ɟ۟ퟘ��#�5�G� �k�}�������^�ׯ �����ʯC�U�g� y���6�����ӿ忐� ���-�?�Q���uχ� �ϫϽ�h������� )���M�_�q߃ߕ�@� �������ߚ��%�7� I�[�������� r������!�3���W� i�{���8��������� ����/ASe �����|� +=�as�� B����/�'/ 9/K/]/o//�/�/�/ �/�/�/�/?#?5?�/ F?k?}?�?�?L?�?�? �?�?O�?1OCOUOgO yO$O�O�O�O�O�O�O 	__-_?_�Oc_u_�_ �_�_V_�_�_�_oo�c�$SMON_�DEFPROG �&���Aa� &*S?YSTEM*obg� $JO0dR�ECALL ?}�Ai ( �}6�copy md:�place_to�rno.tp v�irt:\tem�p\=>10.1�09.25.13:15084 �da4bo�o�o	v}<�e�sumir_barra�o�o�c�ok�}y=�k+sprensa6H[���xxyzrate 61��`���_�q���s8�bfr�s:orderf�il.dat�umpbackE��aV�����}/�db:*.*��ď͏^�p���6t3x��:\&���@8�S�V����}4��a�����eҟc�u��� ����5�P����� ��<�ί_�q�����)� ;�̟ݿ��������J�	�m��w?�fi�ckup*testeir�?ω����� w�o4��K�\�n߀� ��0�B�[����ߑ� �Ǳ���P�a�s� ��3�N�������(� ��L�]�o�����'�9� ʿ�������$ϵ�H� ��k}���+���X ��� ��D��g y����1�T�� ����c/u/�/w }
�11 (/ :/L/�/�/?�&��a �/�/_?q?�?��1 ��?�?O�/�?J 	OmOO���/�ZO �O�O/"/�OF?�Oi_ {_�?�?)O@_V_�_�_ OO�_BO�_eowo
o �O/_�_Ro�o�o_ �o�oP_as��_�_ 3oNo���o(o� Lo]�o����o'9�o �����$��Hڏ k�}���+���X�� ��� ���D�֟g�y�����$SNPX_�ASG 2�������o  0��%����Я  ?���PA�RAM ����� �	��P�Ӥ��Ө$�������OFT_K�B_CFG  �ӣ����OPIN_�SIM  ����}���������R�VNORDY_DOO  )�U����QSTP_DSB�i��ϐ�SR ��� � &�#�D�O�O�:�TO�P_ON_ERR�ʿ��o�PTN ������A���RING_PR�My�ܲVCNT_�GP 2��!���x 	���ϗ��ϰ#��Gߔ�VD��ROP 1��"�8� ��*߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�}�z��� ������������
 C@Rdv��� ���	*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?[?X?j?|? �?�?�?�?�?�?�?!O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo sopo�o�o�o�o�o�o �o 96HZl ~��������� �2�D�V�`�PRG_COUNTJ�s��{�ENB���}�M��L���_UP�D 1'�T  
k�����"�K� F�X�j���������۟ ֟���#��0�B�k� f�x���������ү�� ����C�>�P�b��� ������ӿο��� �(�:�c�^�pςϫ� �ϸ������� ��;� 6�H�Z߃�~ߐߢ��� �������� �2�[� V�h�z�������� ����
�3�.�@�R�{� v������������� *SN`r����t�_INFO� 1�Ҁ� 	 ���3����@�6��3>��>�: ³���A���/^�$C3������BL>?��` @�� Bg���@J� ?&� A-�@9� =�<�Į��4l���A��C�����YSDOEBUG����� �dՉ�SP_PA�SS��B?+L_OG ����  � 9� � �с�UD�1:\;$�<"_M�PCA-셽/�/��x!�/ 쁝&SAV D)��%d!|"��%�(SV�+T�EM_TIME �1D'�� 0�b a^$;�(%  �M7MEMBK  �сd d/�?��?�<X|Ҁ�	 ��9�O:OJLOdmOzI�J
! �;@p1�O�O�O�O�?_@_0_B_T_f_nT�n_ �_�_�_�_�_�_�_o"o\�e1oVohozo�o �o�o�o�o�o�o
 .@Rdv���O5SK�0�8���?�X��F:� 4�HY2OJ�AJ� [@ApJ��A\O����(�O!��Oя���� q��OM�� � �j��@^�p���v_��U����@ӟ���	��� $� C�7og�y��������� ӯ���	��-�?�Q��c�u����������T�1SVGUNSP�D%% '%�T�2MODE_LI�M a9"ܴ2��	� D-۵AS�K_OPTION� �9!F�_DI~ ENB  U��%f�BC2_GRP 2!�u#o2���XB��C����ԼBC?CFG #��*<c #6���`� @I�4�Y��jߣߎ� �߲���������E� 0�i�T��x����� �������/��S�>�w�����t���u��� ��c���	B-f �.��4[ ���� ��� 02D zh������ �/
/@/./d/R/�/ v/�/�/�/�/�(���/ ?&?8?J?�/n?\?~? �?�?�?�?�?�?O�? 4O"OXOFOhOjO|O�O �O�O�O�O�O__._ T_B_x_f_�_�_�_�_ �_�_�_oo>o�/Vo ho�o�o�o(o�o�o�o �o(:Lp^ ��������  �6�$�Z�H�~�l��� ����؏Ə��� �� 0�2�D�z�h���To�� ȟ���
���.��>� d�R�������z�Я�� �����(�*�<�r� `���������޿̿� ��8�&�\�Jπ�n� �ϒϤ������ϴ�� (�F�X�j��ώ�|ߞ� �߲��������0�� T�B�x�f������ ��������>�,�N� t�b������������� ����:(^�v ����H��� $HZl:�~ �������2/  /V/D/z/h/�/�/�/ �/�/�/�/?
?@?.? P?R?d?�?�?�?t�? �?OO*O�?NO<O^O �OrO�O�O�O�O�O�O __8_&_H_J_\_�_ �_�_�_�_�_�_�_o 4o"oXoFo|ojo�o�o �o�o�o�o�o�?6 Hfx���������v&��$T�BCSG_GRP� 2$�u��  �&� 
? ?�  Q�c� M���q��������ˏ���*�1�&8�d�, �F�?&�	� HCA�����b��CS��B�I�����V�>̓�ͪ�n�Ќ�ԝB���333��BElt������AÐ��fff:��.�C����l�?�A���G�w�R���A&� �̧�����@��I� �-���
�X�u�@�R�Р���̻�����	�V3.00I�	'mt7���*� ��%��ֶY��@�ff&� &�H�� qN� �O�  ������ ϏϘ�*�J�21�'8��Ϥ�C�FG )�u�B� E������rd���#��#� I�W��pW�}�hߡߌ� �߰��������
�C� .�g�R��v���� ����	���-��Q�<� u�`�r����������� I�cp"4��g Rw������ 	-?�cN� r��&����� �/</*/`/N/�/r/ �/�/�/�/�/?�/&? ?J?8?Z?\?n?�?�? �?�?�?�?O�? OFO 4OjOXO�O�O`�O�O tO�O_�O0__T_B_ x_f_�_�_�_�_�_�_ �_�_,ooPoboto�o @o�o�o�o�o�o�o�o (L:p^�� ������ �6� $�F�H�Z���~����� ؏Ə����2��OJ� \�n���������� ����
�@�R�d�v� 4���������ί��� �ү(�N�<�r�`��� ������ʿ̿޿�� 8�&�\�Jπ�nϐ϶� ����������"��2� 4�F�|�jߠߎ����� ���� �߼�B�0�f� T��x�������� ����>�,�b�P��� ������v������� :(^L�p� ���� �$ H6lZ|��� ���/�/ /2/ h/�߀/�/�/N/�/�/ �/
?�/.??R?@?v? �?�?�?j?�?�?�?�? O*O<ONOOO�OrO �O�O�O�O�O�O _&_ _J_8_n_\_�_�_�_ �_�_�_�_o�_4o"o XoFoho�o|o�o�o�o �o�o�/$6�/�o xf������ ��,�>���t�b� ������Ώ��򏬏� �&�(�:�p�^����� ����ܟʟ�� �6� $�Z�H�~�l������� دƯ��� ��D�2� T�z�h���Jȿڿ ������
�@�.�d�R� ��vϬϾ����Ϡ�� ����*�`�r߄ߖ� Pߺߨ��������� �&�\�J��n��� ���������"��F� 4�j�X�z�|������� ������0B�Z l~(����� ��,Pbt��D������ s  # &�0/"�$TBJO�P_GRP 2*��� / ?�&	H"O#�,V,����� �� =k% w Ȫ � �� =�$ @ g"	 �CA��&��SC��_%�g!�"G��"k���/�+=�C�S�?��?��&0%0CR  B�4�'??J7�/�/?3�33�2Y&0}?�:;'��v 2�1�0-1E*20�6?�?20��7?C�  D�!�,�� BL��OK:��Z�Bl  @�pB@�� s33C��1 �?gO  A�zG�2jG�&)A)E�OޯJ;��|A?�gff@U@�1C�Z0qzjO�Oz@���U�O�$fff0R)_;^o;xCsQ?ٶ4 )@�O�_tF�X_J\EU<�_�V:�t-�Q(B�*@�Ooh�&-h$o ZGLo6oDoro�o~o8o �o�o�o�o3�o�RlVd��V4��&`�q�%	V3�.00m#mt7A@�s*�l$!�'�� E��qE����E�]\E��HFP=F��{F*HfF�@D�FW�3F�p?F�MF����F�MF���F�şF���F�=F����G�G�.8�CW�R�D3l)D���E"��Ex�
�E��E�,)�FdRFBFH�Fn� F���F��MF�ɽ�F�,
Gl�Gg!G)��G=��GS5��GiĈ;��
�;�o�|& :� @Xz&/��
&"�?�0�&=;-�ESTPARS c (a E#HRw�ABLE 1-V)' @�#R�7�Q � �R�R�R��'#!R�	R�
R��R���!R�R�:R���RDI��`!��ԟ���
�r�Oz���������̯ޮ��Sx�^# <����� ÿտ�����/�A� S�e�wωϛϭϿ��� ����;-w�{�_"��6� �1�C�U���%�7��I�[����NUM [ �`!� �$  ��m���_CFG .���!�@H IMEBF_�TT}���^#��G�V�E10m�H�]�G�R� 1/�� 8$�" �� �A�  ����������� � �2�D�V�h�z��� ����������/
 e@Rhv��� ����*< N`r����� �'///]/8/J/`/�n/�/�/�/�/r���_���t�@~�t�MI__CHANS� ~�� !3DBGLVL�S�~�s�$0ETHERAD ?��w0�"��/�/�?x�?l�$0ROUTq�!�!�4�?�<?SNMASKl8~�>}1255.2E�s�0OBOTO�st�OOL�OFS_DI}���%V9ORQCTRL 0���#��MT�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo&l�OIo8omo�q�PE_DETA�IJ8�JPGL_C�ONFIG 6��ᄀ/ce�ll/$CID$/grp1qo�o�o/壀�?Zl ~���C��� � �2��V�h�z��� ����?�Q����
�� .�@�Ϗd�v������� ��M������*�<� ˟ݟr���������̯@�}a���&�8�J� \���^o��c��`��� ˿ݿ���Z�7�I� [�m�ϑ� ϵ����� �����!߰�E�W�i� {ߍߟ�.��������� ���A�S�e�w�� ���<��������� +���O�a�s������� 8�������'9 ��]o����F ���#5�Y�k}�����`��User V�iew �i}}1�234567890�//,/>/P/X$X� �cx/���2� U�/�/�/�/??s/�/�3�/b?t?�?�? �?�??�?�.4Q?O (O:OLO^OpO�?�O�.5O�O�O�O __$_�OE_�.6�O~_�_�_@�_�_�_7_�_�.7m_ 2oDoVohozo�o�_�o�.8!o�o�o
.�@�oagr l�Camera ��o����� �ޢE�*�<�N��h��z��������I   �v�)��$�6�H�Z� l����������؟� ��� �2�Y��vP9 ɟ~�������Ưد� ��� �k�D�V�h�z� ����E�W�I5���� � �2�D��h�zό� ׿����������
߱� W�ދ��X�j�|ߎߠ� ��Y�������E��0� B�T�f�x�߁ulY� ��������
����@� R�d������������ ����W� iy�.@R dv�/���� �*<N��W� �i������� �/*/</�`/r/�/ �/�/�/as9F/�/ ??1?C?U?�f?�? �?D/�?�?�?�?	OO-O�j	�u0�?hOzO �O�O�O�Oi?�O�O
_ �?._@_R_d_v_�_/O AO�p�{,_�_�_oo )o;o�O_oqo�o�_�o �o�o�o�o�_�u�� �oM_q���No ���:�%�7�I� [�m�NEa����ˏ ݏ����7�I�[� ���������ǟٟ�� ��ͻp�%�7�I�[�m� �&�����ǯ���� �!�3�E�쟒�9�ܯ ������ǿٿ뿒�� !�3�~�W�i�{ύϟ� ��X�����H����!� 3�E�W���{ߍߟ��π������������  ��L�^�p�� ���������� ��   "�*�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/�</N/`/r/�/�  }
��(  �@�( 	 �/�/�/ �/�/? ?6?$?F?H?�Z?�?~?�?�?�?�*2� �l�O/OAO ��eOwO�O�O�O�O�� O�O�O_TO1_C_U_ g_y_�_�O�_�_�__ �_	oo-o?oQo�_uo �o�o�_�o�o�o�o ^opoM_q�o� �����6�%� 7�~[�m�������� �ُ���D�!�3�E� W�i�{�ԏ��ß՟ �����/�A�S��� w�����⟿�ѯ��� ��`�=�O�a����� ������Ϳ߿&�8�� '�9π�]�oρϓϥ� ����������F�#�5� G�Y�k�}��ϡ߳��� �������1�C�� ��y����������� ��	��b�?�Q�c��� ������������(� )p�M_q��8����0@ �������� ���#frh:\tp�gl\robots\m10ia4_7l.xml� Xj|�������.��/1/C/ U/g/y/�/�/�/�/�/ �/�//?-???Q?c? u?�?�?�?�?�?�?�? 
?O)O;OMO_OqO�O �O�O�O�O�O�OO _ %_7_I_[_m__�_�_ �_�_�_�__�_!o3o EoWoio{o�o�o�o�o �o�o�_�o/AS ew������ �o��+�=�O�a�s� ��������͏ߏ��I �<�<  ?� �4��,�N�|�b��� ����ʟ�Ο���0� �8�f�L�~�������趯�����(�$�TPGL_OUT?PUT 9����w� $� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ������$����2345?678901���  �2�D�V�^����υ� �ߩ߻�����w���� '�9�K�]���}g�� �������o���� 1�C�U�g���u����� ������}���-? Qc������ ���);M_ q	����� ��%/7/I/[/m// /�/�/�/�/�/�/�/ ?3?E?W?i?{??%? �?�?�?�?�?O�?O AOSOeOwO�O!O�O�O��O�O�O_�O� $$Ӣ��OW=_ o_a_�_�_�_�_�_�_ �_�_#ooGo9oko]o �o�o�o�o�o�o�o�o C5g}��@������}@���"�� ( 	 iW�E�{�i��� ��Ï��ӏՏ��� A�/�e�S���w����� ���џ���+��;��=�O���s����Ƹ ? <<\ޯ �)�ͯ�)��M�_� ��ʯ����<���ؿ�� Ŀ� �~�$�V��B� �Ϟ�x�����2ϼ�
� ����@�R�,�v߈��� p߾���j������� <�߬�r����� ������`�&�8��� $�n�H�Z�������� ������"4Xj ��R��L��� �|Tf � �v��0B// �&/P/*/</�/�/� �/�/h/�/??�/:? L?�/4?�??n?�?�? �?�? O^?�?6OHO�? lO~OXO�O�OO$O�O �O�O_2___h_z_ �O�_�_J_�_�_�_�_�o.o��)WGL�1.XML�cm��$TPOFF_L�IM Š�p����qfN_SV�y`  �t�jP_MON :��S�d�p�p2mi�STRTCHK �;���f~tbVTCOMPAT�h�*q�fVWVAR �<�mMx�d � e�p�b�ua_DEFPRO�G %�i%�SEGURA_B�AR�pRECEP�TOR�rISP�LAY�`�n�rIN�ST_MSK  ��| �zINU�SE�p"�rLCK�)��{QUICKM�ENM��tSCRE�l���+rtpsc�t)������b���_��STz�iR�ACE_CFG �=�iMt�`	�nt
?��HNL� 2>�z���T{  zr@�R�d�v����������К�ITEM �2?,� �%$�12345678�90�%�  =<��C�U�]�  !c�k�wp'���ns� ѯ5����k������ j�ů��鯕���A�1� C�U�o�y�󿝿I�o� ��忥�	��-ϧ�Q� ��#�5ߙ�A߽����� e߳������M���q� ��L��g��ߋ��� ��%�w� �[���+� Q�c���o�������� 3���{�;���� ��G_����/� Se.�I�m ���=�a /3/������ k//�/�/�/]/?�/ �/�/?�/u?�?�?? �?5?G?Y?�?+O�?OO aO�?mO�?�?�OO�O CO__yO+_�O�Ox_ �O�_�O�_�_�_?_�_ c_u_�_o�_Wo}o�o �_�oo)o;o�o�oqo 1C�oO�o�o� �%��[���Z��S�@��_�ψ  ے_� 8����y
 Ï��Џ���UD1:�\���q�R_G�RP 1A �?� 	 @�pe� w�a���������ߟ͞����ّ�>�)�<b�M�?�  }��� y�����ӯ������ 	��Q�?�u�c�����0����Ϳ�	-����o�SCB 2B{� h�e�wωπ�ϭϿ�������e�U�TORIAL �C{��@�j�V_C�ONFIG D�{���������O�OUTPUT E{���������� �%�7�I�[�m��� ������������ %�7�I�[�m������ ����������!3 EWi{���� ����/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/��/? ?'?9?K?]?o?�?�? �?�?�?�/�?�?O#O 5OGOYOkO}O�O�O�O �O�O�?�O__1_C_ U_g_y_�_�_�_�_�_ �O�_	oo-o?oQoco uo�o�o�o�o�o�_�o );M_q� �����yߋ��� �-�?�Q�c�u����� ����Ϗ���o�)� ;�M�_�q��������� ˟ݟ� ��%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� 
��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ���1CUgy �������	 -?Qcu��������/�x���$/6/ !/ a/��/�/�/�/�/�/ �/??'?9?K?]? �?�?�?�?�?�?�?�? O#O5OGOYOkO|?�O �O�O�O�O�O�O__ 1_C_U_g_xO�_�_�_ �_�_�_�_	oo-o?o Qocot_�o�o�o�o�o �o�o);M_ q�o������ ��%�7�I�[�m�~ ������Ǐُ���� !�3�E�W�i�z����� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o��~��$TX_SCREEN 1F8%�  �}�~���������
����m&��\�n߀ߒ� �߶�-�?������"� 4�F��j��ߎ��� ������_����0�B� T�f�x��������� ������>��b t����3�W (:L^�� ������e/ �6/H/Z/l/~/�//��/�$UALRM_MSG ?����� �/���/�/ )??M?@?q?d?v?�?��?�?�?�?�?O�%S�EV  �-�EF�"ECFG �H����  ���@�  AuA �  Bȁ�
  O���ŨO�O�O�O�O __&_8_J_\_jWQA�GRP 2I[K; 0��	 �O�_�� I_BBL_N�OTE J[JT��l������g@�RDEF�PRO� %�+ �(%MAIN �A_PRENSA VISION�_%OVoAozoeo�o�o �o�o�o�o�o@��[FKEYDAT�A 1K�ɞPp jG���_��0����z,(�����([ INS�T ]'�)�  I�RECTS�~��N�Dh���b�ES I�CEB���[ED�CMDƏ��ORE<�FO��C�U� <�y�`�������ӟ�����	��-��Q�c�� ��/frh�/gui/whi�tehome.pngd�����Ưد�{�{�inst����/�A�S�e���  >|�direc����������п�q���in���.�@�R�d�v���yes��ϲϰ�������π{�edcmd��#�5�G߸Y�k�}� �{�arwrgϲ����� ���߁��)�;�M�_� q����������� ���%�7�I�[�m�� ������������� ��3EWi{� ������/ ASew��r�� ����/!/(E/ W/i/{/�/�/./�/�/ �/�/??�//?S?e? w?�?�?�?<?�?�?�? OO+O�?OOaOsO�O �O�O8O�O�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o �_Goko}o�o�o�o�o To�o�o1C�o gy����P� �	��-�?�Q��u�@��������Ϗj�܋�u�܏�(�s��Q�c�r�,I���A��POINT M|����  OOKß��G�AREL  �T�� CHOI�CE]��TOUCHUPG�H�s� ��~�����߯�د� ��9�K�2�o�V�����茿ɿ��whi?tehome���� �2�D�V�	�poin�ߍϟϱ�����`��look}����(�:�L�^���pgkarel}Ϙߪ߼��������choic ���� �2�D�V�h�k���touchup�ߠ��������g�}�arwrg|� "�4�F�X�j�a����� ��������w�0 BTfx��� ����,>P bt����� �/�(/:/L/^/p/ �//�/�/�/�/�/ ? ׿�/6?H?Z?l?~?�? �/�?�?�?�?�?O�? 2ODOVOhOzO�O�O-O �O�O�O�O
__�O@_ R_d_v_�_�_)_�_�_ �_�_oo*o�_No`o ro�o�o�o7o�o�o�o &�oJ\n� ���E���� "�4��X�j�|����� ��A�֏�����0� B�яf�x��������� O������,�>�ټ�L������u�����q���ͯ��,������"�	�F� X�?�|�c�������ֿ ������0��T�f� Mϊ�qϮϕ������� ���,�>�?b�t߆� �ߪ߼�˟������ (�:�L���p���� ����Y��� ��$�6� H���l�~��������� ��g��� 2DV ��z�����c �
.@Rd� ������q/ /*/</N/`/��/�/ �/�/�/�/�//?&? 8?J?\?n?�/�?�?�? �?�?�?{?O"O4OFO XOjO|OSߠO�O�O�O �O�OO_0_B_T_f_ x_�__�_�_�_�_�_ o�_,o>oPoboto�o o�o�o�o�o�o �o:L^p��# ���� ���6� H�Z�l�~�����1�Ə ؏���� ���D�V� h�z�����-�ԟ� ��
��.���R�d�v� ������;�Я���� �*���N�`�r�����h�����@����@������	��+�=��,)�n�!� ��y϶��ϯ������ "�	�F�-�j�|�cߠ� �����߽������� B�T�;�x�_���O ��������,�;�P� b�t���������K��� ��(:��^p ����G��  $6H�l~� ���U��/ / 2/D/�h/z/�/�/�/ �/�/c/�/
??.?@? R?�/v?�?�?�?�?�? _?�?OO*O<ONO`O �?�O�O�O�O�O�OmO __&_8_J_\_�O�_ �_�_�_�_�_�_��o "o4oFoXojoq_�o�o �o�o�o�o�o�o0 BTfx��� �����,�>�P� b�t��������Ώ�� ����(�:�L�^�p� �������ʟܟ� � ���6�H�Z�l�~��� ���Ưد������ 2�D�V�h�z�����-� ¿Կ���
�ϫ�@� R�d�vψϚ�)Ͼ���@������*�`,���`����U�g�y�Qߛ߭߇�, ���ߑ����&�8�� \�C���y����� �������4�F�-�j� Q���u����������� �_BTfx� ������� ,�Pbt��� 9���//(/� L/^/p/�/�/�/�/G/ �/�/ ??$?6?�/Z? l?~?�?�?�?C?�?�? �?O O2ODO�?hOzO �O�O�O�OQO�O�O
_ _._@_�Od_v_�_�_ �_�_�___�_oo*o <oNo�_ro�o�o�o�o �o[o�o&8J \3������ �o��"�4�F�X�j� �������ď֏�w� ��0�B�T�f����� ������ҟ������ ,�>�P�b�t������ ��ί�򯁯�(�:� L�^�p��������ʿ ܿ� Ϗ�$�6�H�Z� l�~�Ϣϴ������� ��ߝ�2�D�V�h�z� ��߰���������
� ��.�@�R�d�v����qp���qp���������������,	N�r�Y� �������������� &J\C�g� ������"4 X?|�m�� ���/�0/B/T/ f/x/�/�/+/�/�/�/ �/??�/>?P?b?t? �?�?'?�?�?�?�?O O(O�?LO^OpO�O�O �O5O�O�O�O __$_ �OH_Z_l_~_�_�_�_ C_�_�_�_o o2o�_ Vohozo�o�o�o?o�o �o�o
.@�od v����M�� ��*�<��`�r��� ������̏����� &�8�J�Q�n������� ��ȟڟi����"�4� F�X��|�������į ֯e�����0�B�T� f�����������ҿ� s���,�>�P�b�� �ϘϪϼ������ρ� �(�:�L�^�p��ϔ� �߸�������}��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z�	��������������
��>����5G Y1{�g,y� q���<# `rY�}��� ��/&//J/1/n/ U/�/�/�/�/�/�/�/ ݏ"?4?F?X?j?|?�� �?�?�?�?�?�?O�? 0OBOTOfOxO�OO�O �O�O�O�O_�O,_>_ P_b_t_�_�_'_�_�_ �_�_oo�_:oLo^o po�o�o#o�o�o�o�o  $�oHZl~ ��1�����  ��D�V�h�z����� ��?�ԏ���
��.� ��R�d�v�������;� П�����*�<�? `�r�����������ޯ ���&�8�J�ٯn� ��������ȿW���� �"�4�F�տj�|ώ� �ϲ�����e����� 0�B�T���xߊߜ߮� ����a�����,�>� P�b��߆������ ��o���(�:�L�^� ��������������� }�$6HZl�� ������y� 2DVhzQ��|�Q�����������,�/./�/R/9/v/�/ o/�/�/�/�/�/?�/ *?<?#?`?G?�?�?}? �?�?�?�?OO�?8O O\OnOM��O�O�O�O �O�O�_"_4_F_X_ j_|__�_�_�_�_�_ �_�_o0oBoTofoxo o�o�o�o�o�o�o �o,>Pbt� �������(� :�L�^�p�����#��� ʏ܏� ����6�H� Z�l�~������Ɵ؟ ���� ���D�V�h� z�����-�¯ԯ��� 
����@�R�d�v��� �����Oп����� *�1�N�`�rτϖϨ� ��I�������&�8� ��\�n߀ߒߤ߶�E� �������"�4�F��� j�|������S��� ����0�B���f�x� ����������a��� ,>P��t�� ���]�( :L^����� ��k //$/6/H/ Z/�~/�/�/�/�/�/��/���+������?'?9=?[?m?G6,YO�?QO�? �?�?�?�?OO@ORO 9OvO]O�O�O�O�O�O �O_�O*__N_5_r_ �_k_�_�_�_�_��o o&o8oJo\ok/�o�o �o�o�o�o�o{o" 4FXj�o��� ���w��0�B� T�f�x��������ҏ ������,�>�P�b� t��������Ο��� ���(�:�L�^�p��� �����ʯܯ� ��� $�6�H�Z�l�~���� ��ƿؿ���ϝ�2� D�V�h�zό�ϰ��� ������
���_@�R� d�v߈ߚߡϾ����� ����*��N�`�r� ����7�������� �&���J�\�n����� ����E�������" 4��Xj|��� A���0B �fx����O ��//,/>/�b/ t/�/�/�/�/�/]/�/ ??(?:?L?�/p?�? �?�?�?�?Y?�? OO�$O6OHOZO�$UI�_INUSER � ���{A��  �[O_O_MENHI�ST 1L{E�  ( ��@��'/SO�FTPART/G�ENLINK?c�urrent=m�enupage,98,1�O__0_�B_ �7�O�Eed�it�BCOLOC�A_BARRA_TORNO�O�_�_��_�32X_j_|SPRENSA�_o/oAo�8�O�O71`o�o��o�o�o�;`o�^S�EGU�P�SRECEP�P,1�o/A�S�9�o�_|USE�_IRVISIOANo����1)hz~MAI�#�5�G��Y��0(��N148�,2\�����͏ߏ���0�A����"�4�F�X�j� �������� şן�x���1�C� U�g�����������ӯ ������-�?�Q�c� u��������Ͽ�� ���)�;�M�_�qσ� ϧϹ��������� %�7�I�[�m�ߑߔ� ������������3� E�W�i�{������ ����������A�S� e�w�����*������� ����=Oas ���8��� '�0]o�� ������/#/ 5/�Y/k/}/�/�/�/ B/�/�/�/??1?C? �/g?y?�?�?�?�?P? �?�?	OO-O?O�?PO uO�O�O�O�O�O^O�O __)_;_M_8�O�_ �_�_�_�_�_�Ooo %o7oIo[o�_o�o�o �o�o�o�ozo!3 EWi�o���� ��v��/�A�S� e�w��������я� �����+�=�O�a�s��^[�$UI_PA�NEDATA 1�N������  	�}�c/frh/cg�tp/flexd�ev.stm?_�width=0&�_height=�10ԐŐice=�TP&_line�s=3Ԑcolu�mns=4Ԑfo�nܐ4&_pag�e=doubŐ1���\V)prim#�L�  }O�s���0������ͯ )ϯ� گ���;�M�4�q�X� ������˿������%�\V�� �E�eP�1�]�d���ɟ۞2����2</�-�dual���� _��"�4�F�X�j�� ��u߲��߫������ ��B�)�f�M���؃���3� G�2T �����*�<�N�`� ����Ϩ��������� i�&8\C� �y�����@�4Xj=� �� ����������  /S$/��H/Z/l/~/ �/�/	/�/�/�/�/�/  ?2??V?=?z?a?�? �?�?�?�?�?
O}� @OROdOvO�O�O�?�O 1/�O�O__*_<_N_ �Or_Y_�_}_�_�_�_ �_�_o&ooJo1ono �ogo�oO)O�o�o�o "4�oXj�O� �����O�� 0�B�)�f�M������� �������ݏ��>� �o�o���������Ο ��3��w(�:�L�^� p���韦�����ܯï  ����6��Z�A�~� ��w�����ؿ�]�o�  �2�D�V�h�z�Ϳ�� ���������
��.� ��R�9�v�]ߚ߬ߓ� �߷������*��N� `�G����	������ �������"�)��G� ��6�s����������� 4�������K2 oV���������#�����$�UI_POSTY�PE  �� 	 /��UQUICKM_EN  ds��WRESTOR�E 1O�  �B�� /#���m+/ T/f/x/�/�/?/�/�/ �/�/?�/,?>?P?b? t?/�?�?�??�?�? OO(O�?LO^OpO�O �O�OIO�O�O�O __ �?_1_C_�O~_�_�_ �_�_i_�_�_o o2o �_Vohozo�o�oI_So �o�oAo�o.@R d�����s ���*�<��oI�[� m������̏ޏ���� �&�8�J�\�n����ट��ȟڟ�SCR�E�?��u1sc�u2��3�4�5�6��7�8��TAT`� ��M�USER�����k�s���3��4��5*��6��7��8��U�NDO_CFG �Pd����UPD�X����N�one���_IN_FO 1Q�<��0%��W���E� ��i���������տ ���:�L�/�pς�e���ύ)�OFFSEOT Td@��� {������	��-�Z� Q�cߐ߇ߙ��ϝ��� ���� ��)�V�M�_�@q�۹�����
����t��)�WORK U4�����A��S��ψ�UFRAM�E  ���&�R�TOL_ABRT8��$���ENB����?GRP 1V��Cz  A� ��+=Oas�����U������?MSK  �<����N��%4��%x��)��_EVN��b���>�2W���
 h��UE�V��!td:\�event_usger\-�C7�d��}�F��SP���spotwe{ld�!C6����!�Z/ �/:'�H/~/l/�/�/ �/�/-?�/Q?�/? ? �?D?�?h?z?�?O�? )O�?�?OqO`O�O@O RO�OvO�O_�O�O7_��O[__Z]W+�2X����8V_�_�_ �_�_o�_,o>oo botoOo�o�o�o�o�o �o�o:L'p��]����$V�ARS_CONFuI�Y�� FP{�{��|CCRG�C\��>�{�t�]D� BH� pk��a�C�� ��}�?񀏀C,&Q=��Ͷ��A �MR2�b���	}�	���@�%1: S�C130EF2 Q*����{�����X�� �5}�����A�@k�C�F� w�Q�[���|����������T����\��ϟ �\� B���;�e�@�ǟ`� ����S�����̯��� ۯ�&�}��\�G�Y����E���ȿ�TCC��c
���������pGF�pgd���-�23456789017�?��ׁ$���4�v�Nm�� ��϶�BW������i�}�:�o=L A�څ�6�@�6�ͿZ�H��i�7����(��W� ��-�]�X�jĈߚߕ� �Ϲ���������%� 7�I�r�m�ߨ�ߵ� ���������8�3�E� W������}������� ������/�A�S�e�<w��MODE��t� �RSLT 3e�|k�%"zς� �;�1��d��`|��SELEC���c��	IA_W�O�Pf ��� W,		�������G�P ������RTSYN'CSE� ��$�	#�WINURL ?*ـ�;\/n/��/�/�/�/�uISI?ONTMOU����A# ��%�gSۣ�SۥP�� FR:\�#�\DATA\�/ �� MC6�LOG?   7UD16EX@?\��' B@ ���2T1���?T1�?��?����� n?6  ���GV�2�\� -��5��   ��Z�@U0}58TRAINj?h��*B{Rd_Cp��NF#`{2�'$t�"��h#� (� kI�Mw��O�O�O�O�O 1__U_C_]_g_y_�_��_�_�(STA� i���@�?o0oI:$�obo�%_GE�jv#��~@ �
��\��btgHOMIN��kSۮ��`�P2,,��CWǖB�veJMPERR {2l#�
  Qo I:��"�4Fwj |����������&%S_g0REr�m�^۴LEXd�n�1-ehoV�MPHASE  ��e׃BޱOF�F _ENB  ��$VP2�$o/Sۯ��x�c C;�@ �@�;����?s33'D*AA ��]� ��0ޱ�`r}�XC��܅���p\A-۟E �� ����#�5������� ������}�������� ��c�X���A����� ϯ�+��߿��M� B�q���xϊϹ���� ��������7�I�;�m� b�)ߣ�Eߓߡ߳��� ��3���W�L�{ߍ� �ߑ���������� /�$�6�e�W���c�y� ������������� O���?M_q��� ����'9�= 7Is����� �/m/%/3/E/�s�TD_FILTuE�`s�k �x2�`����/�/�/�/ �/	??-???Q?�6�/ ~?�?�?�?�?�?�?�?�O OoiSHIFTMENU 1t}<5�%5�~O)�\O �O�O�O�O�O�O�O'_ �O_6_o_F_X_�_|_��_�_�_	LIV�E/SNAP�S?vsfliv���_��z`ION �ҀU
`bmenu &o+o�_�o�oV"<E�uz��4IMO�v����zq�WAIT�DINEND  a�ec��b�fOKوNOUT�hSD�yTIMdu��o|G�}#�{C�z�b�z�xRELE���ڋxTM�{�d=��c_ACT`و���x_DATA �wz���%  E�GA_TORNOx�o.Mx�RDIS
`~E��$XVR�a�x�n�$ZAB�C_GRP 1yvz��� ,��2̏.MZD��CSKCH�`z���aP@��h@�IP�b{'���şן�[��MPCF_G 1|'���0�r�8�d�� �}'��p�s�� 	(���  �<l0  �F���>�:X��L"?!h>���h�3���͋�M��5<=�<�Į��4l�>�w����?��C�=@H����! ?c�"������ɯۯ���?��o���w����� /����A��C�˿ݸĸ����	��P1�?�i��[�#���l����<'��+�?=�B�=ĺ������0?��?4��E�D�!@H�����?c#ײX�	��`~����_CYLIND~!�� Р ,(  *.�?ݧ`+�h�Oߌ�s� �� ������(�	�x�-�� &�c�߇������� j�P����)��~�_��q��� �2�'��� �&�����������&��I��cA����SPHERE 2������ ����A�T/A ��e����� �/N`=/�a/ H/Z/�/��/�/�/�ZZ� ��f